-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity OndraViLi_v27 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(11 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of OndraViLi_v27 is


  type ROM_ARRAY is array(0 to 4095) of std_logic_vector(7 downto 0);
  constant ROM : ROM_ARRAY := (
    x"F3",x"31",x"90",x"D4",x"C3",x"CD",x"18",x"E9", -- 0x0000
    x"E1",x"22",x"E3",x"D4",x"C9",x"30",x"32",x"37", -- 0x0008
    x"C3",x"A0",x"D4",x"25",x"F8",x"C3",x"33",x"1D", -- 0x0010
    x"E3",x"F5",x"7E",x"23",x"D7",x"F1",x"E3",x"C9", -- 0x0018
    x"DF",x"01",x"7C",x"D7",x"DF",x"02",x"18",x"2A", -- 0x0020
    x"E5",x"D5",x"ED",x"5B",x"38",x"D6",x"18",x"25", -- 0x0028
    x"7C",x"87",x"67",x"87",x"D6",x"F9",x"18",x"26", -- 0x0030
    x"E5",x"D5",x"C5",x"F5",x"CD",x"B5",x"D5",x"CD", -- 0x0038
    x"A4",x"18",x"CD",x"C9",x"1A",x"3A",x"27",x"D6", -- 0x0040
    x"CB",x"8F",x"D3",x"03",x"F1",x"C1",x"D1",x"E1", -- 0x0048
    x"FB",x"C9",x"7D",x"D7",x"C9",x"19",x"CD",x"4F", -- 0x0050
    x"1F",x"7E",x"B7",x"D1",x"E1",x"C9",x"84",x"2F", -- 0x0058
    x"65",x"6F",x"7C",x"2F",x"67",x"C9",x"CD",x"CD", -- 0x0060
    x"D5",x"ED",x"7B",x"C2",x"D4",x"21",x"00",x"00", -- 0x0068
    x"22",x"0A",x"D6",x"22",x"08",x"D6",x"3E",x"0F", -- 0x0070
    x"32",x"28",x"D6",x"3E",x"04",x"D3",x"03",x"3A", -- 0x0078
    x"08",x"E0",x"4F",x"AF",x"D3",x"03",x"32",x"27", -- 0x0080
    x"D6",x"CB",x"51",x"28",x"40",x"ED",x"56",x"FB", -- 0x0088
    x"CB",x"61",x"2A",x"02",x"D6",x"28",x"0A",x"CB", -- 0x0090
    x"49",x"2A",x"9E",x"D5",x"28",x"03",x"2A",x"04", -- 0x0098
    x"D6",x"C3",x"E5",x"D4",x"21",x"2F",x"D6",x"34", -- 0x00A0
    x"23",x"35",x"F0",x"36",x"00",x"EB",x"21",x"2E", -- 0x00A8
    x"D6",x"7E",x"E6",x"06",x"FE",x"02",x"C0",x"3A", -- 0x00B0
    x"E0",x"D4",x"12",x"3A",x"27",x"D6",x"E6",x"F9", -- 0x00B8
    x"D3",x"03",x"ED",x"5B",x"36",x"D6",x"2A",x"38", -- 0x00C0
    x"D6",x"19",x"C3",x"AF",x"D4",x"3E",x"6B",x"D3", -- 0x00C8
    x"0A",x"3E",x"30",x"D3",x"03",x"3E",x"14",x"DB", -- 0x00D0
    x"09",x"3E",x"7A",x"DB",x"3D",x"3E",x"B2",x"DB", -- 0x00D8
    x"5A",x"3E",x"10",x"D3",x"03",x"3E",x"2F",x"DB", -- 0x00E0
    x"08",x"AF",x"DB",x"80",x"3E",x"20",x"D3",x"03", -- 0x00E8
    x"3E",x"29",x"DB",x"1C",x"AF",x"DB",x"80",x"21", -- 0x00F0
    x"A0",x"D5",x"E5",x"AF",x"77",x"23",x"BC",x"20", -- 0x00F8
    x"FB",x"E1",x"06",x"20",x"36",x"C9",x"23",x"23", -- 0x0100
    x"23",x"10",x"F9",x"21",x"BF",x"19",x"11",x"A0", -- 0x0108
    x"D4",x"01",x"DE",x"00",x"ED",x"B0",x"21",x"9D", -- 0x0110
    x"1A",x"06",x"05",x"5E",x"23",x"51",x"EB",x"3E", -- 0x0118
    x"C3",x"CD",x"18",x"D5",x"1A",x"13",x"23",x"CD", -- 0x0120
    x"18",x"D5",x"1A",x"13",x"23",x"CD",x"18",x"D5", -- 0x0128
    x"EB",x"10",x"E8",x"CD",x"C3",x"1E",x"21",x"41", -- 0x0130
    x"19",x"06",x"19",x"CD",x"CE",x"22",x"C3",x"69", -- 0x0138
    x"18",x"1F",x"03",x"02",x"0B",x"20",x"5A",x"64", -- 0x0140
    x"72",x"61",x"76",x"C9",x"20",x"56",x"C1",x"73", -- 0x0148
    x"20",x"4F",x"4E",x"44",x"52",x"41",x"20",x"04", -- 0x0150
    x"0D",x"0D",x"DF",x"0D",x"01",x"5C",x"19",x"C5", -- 0x0158
    x"DF",x"1B",x"DF",x"46",x"2A",x"BE",x"D4",x"CD", -- 0x0160
    x"DD",x"23",x"11",x"32",x"D5",x"06",x"00",x"CD", -- 0x0168
    x"CE",x"20",x"CD",x"9E",x"21",x"20",x"1E",x"57", -- 0x0170
    x"CD",x"8C",x"19",x"6F",x"CD",x"8C",x"19",x"67", -- 0x0178
    x"15",x"28",x"15",x"15",x"20",x"0B",x"CD",x"D6", -- 0x0180
    x"22",x"C3",x"E5",x"D4",x"CD",x"9E",x"21",x"C8", -- 0x0188
    x"F1",x"DF",x"3F",x"DF",x"0D",x"C3",x"D6",x"22", -- 0x0190
    x"CD",x"8C",x"19",x"4F",x"CD",x"8C",x"19",x"47", -- 0x0198
    x"CD",x"8C",x"19",x"CD",x"18",x"D5",x"ED",x"A1", -- 0x01A0
    x"EA",x"A0",x"19",x"18",x"C5",x"01",x"80",x"0A", -- 0x01A8
    x"21",x"28",x"D6",x"7E",x"E6",x"1F",x"B1",x"77", -- 0x01B0
    x"FB",x"76",x"10",x"FD",x"A9",x"77",x"C9",x"C3", -- 0x01B8
    x"CD",x"1C",x"C3",x"62",x"1F",x"C3",x"AB",x"1F", -- 0x01C0
    x"C3",x"85",x"20",x"C3",x"50",x"20",x"C3",x"3B", -- 0x01C8
    x"20",x"C3",x"78",x"1E",x"C3",x"69",x"18",x"69", -- 0x01D0
    x"00",x"57",x"CC",x"58",x"CC",x"A0",x"CF",x"A0", -- 0x01D8
    x"D3",x"A0",x"D4",x"6B",x"1F",x"13",x"0C",x"0B", -- 0x01E0
    x"0B",x"00",x"1F",x"00",x"16",x"00",x"0F",x"00", -- 0x01E8
    x"1F",x"00",x"1F",x"00",x"00",x"00",x"01",x"00", -- 0x01F0
    x"0F",x"00",x"1F",x"00",x"1F",x"02",x"19",x"19", -- 0x01F8
    x"28",x"15",x"F6",x"1C",x"CD",x"E9",x"D4",x"E9", -- 0x0200
    x"E5",x"21",x"27",x"D6",x"CB",x"CE",x"F5",x"7E", -- 0x0208
    x"D3",x"03",x"F1",x"E1",x"C9",x"ED",x"53",x"06", -- 0x0210
    x"D6",x"E3",x"5E",x"23",x"56",x"23",x"E3",x"E5", -- 0x0218
    x"21",x"E9",x"D4",x"E3",x"D5",x"ED",x"5B",x"06", -- 0x0220
    x"D6",x"E5",x"21",x"27",x"D6",x"CB",x"8E",x"18", -- 0x0228
    x"DD",x"CD",x"E9",x"D4",x"7E",x"18",x"F2",x"CD", -- 0x0230
    x"E9",x"D4",x"77",x"18",x"EC",x"F5",x"AF",x"D3", -- 0x0238
    x"03",x"FF",x"3A",x"27",x"D6",x"CB",x"CF",x"D3", -- 0x0240
    x"03",x"F1",x"C9",x"E7",x"66",x"18",x"C9",x"CF", -- 0x0248
    x"10",x"4B",x"EF",x"44",x"E3",x"F5",x"7E",x"23", -- 0x0250
    x"FE",x"12",x"38",x"04",x"F1",x"E3",x"18",x"71", -- 0x0258
    x"E5",x"D5",x"5F",x"16",x"00",x"21",x"5A",x"D5", -- 0x0260
    x"19",x"19",x"7E",x"23",x"66",x"6F",x"22",x"57", -- 0x0268
    x"D5",x"D1",x"E1",x"F1",x"E3",x"E7",x"00",x"00", -- 0x0270
    x"C9",x"10",x"18",x"BE",x"D5",x"BD",x"1A",x"AC", -- 0x0278
    x"1A",x"44",x"1C",x"1E",x"24",x"DD",x"23",x"B0", -- 0x0280
    x"19",x"CE",x"20",x"32",x"22",x"9E",x"21",x"5C", -- 0x0288
    x"22",x"E2",x"22",x"D6",x"22",x"C2",x"1B",x"C3", -- 0x0290
    x"1E",x"5A",x"19",x"28",x"18",x"38",x"1E",x"D5", -- 0x0298
    x"20",x"F6",x"D4",x"00",x"30",x"D5",x"08",x"35", -- 0x02A0
    x"D5",x"66",x"2C",x"D5",x"E5",x"C5",x"21",x"27", -- 0x02A8
    x"D6",x"4E",x"CB",x"C6",x"CD",x"BD",x"1A",x"28", -- 0x02B0
    x"FB",x"71",x"C1",x"E1",x"C9",x"E5",x"D5",x"C5", -- 0x02B8
    x"FB",x"CD",x"5E",x"1B",x"B7",x"C1",x"D1",x"E1", -- 0x02C0
    x"C9",x"3A",x"28",x"D6",x"D3",x"0A",x"3A",x"27", -- 0x02C8
    x"D6",x"CB",x"D7",x"CB",x"8F",x"D3",x"03",x"21", -- 0x02D0
    x"01",x"E0",x"7E",x"E6",x"0B",x"CC",x"B5",x"D4", -- 0x02D8
    x"2E",x"05",x"7E",x"E6",x"07",x"CC",x"BB",x"D5", -- 0x02E0
    x"21",x"1D",x"D6",x"7E",x"B7",x"28",x"01",x"35", -- 0x02E8
    x"3A",x"09",x"D6",x"F5",x"B7",x"C4",x"A0",x"D5", -- 0x02F0
    x"F1",x"E6",x"10",x"C0",x"21",x"1C",x"D6",x"35", -- 0x02F8
    x"F0",x"34",x"21",x"CA",x"D4",x"11",x"09",x"E0", -- 0x0300
    x"1A",x"E6",x"1F",x"47",x"A6",x"0E",x"80",x"20", -- 0x0308
    x"0F",x"78",x"B6",x"EE",x"1F",x"0E",x"00",x"20", -- 0x0310
    x"07",x"23",x"23",x"1D",x"F2",x"08",x"1B",x"C9", -- 0x0318
    x"16",x"80",x"CB",x"02",x"0C",x"0F",x"30",x"FA", -- 0x0320
    x"7A",x"AE",x"77",x"23",x"7A",x"A6",x"20",x"02", -- 0x0328
    x"CB",x"F1",x"7B",x"87",x"87",x"83",x"81",x"4F", -- 0x0330
    x"21",x"09",x"D6",x"34",x"23",x"CD",x"51",x"1B", -- 0x0338
    x"71",x"3E",x"02",x"32",x"1C",x"D6",x"CB",x"79", -- 0x0340
    x"C0",x"3A",x"28",x"D6",x"F6",x"E0",x"D3",x"0A", -- 0x0348
    x"C9",x"7E",x"3C",x"E6",x"0F",x"77",x"6F",x"26", -- 0x0350
    x"00",x"11",x"0C",x"D6",x"19",x"C9",x"CD",x"D3", -- 0x0358
    x"D5",x"CD",x"44",x"1C",x"21",x"1D",x"D6",x"20", -- 0x0360
    x"18",x"7E",x"B7",x"3E",x"00",x"C0",x"3A",x"08", -- 0x0368
    x"D6",x"07",x"3E",x"00",x"D0",x"3A",x"28",x"D6", -- 0x0370
    x"F6",x"E0",x"D3",x"0A",x"3A",x"DE",x"D4",x"18", -- 0x0378
    x"0C",x"CB",x"77",x"C2",x"11",x"1C",x"2F",x"32", -- 0x0380
    x"08",x"D6",x"3A",x"DF",x"D4",x"77",x"CD",x"A1", -- 0x0388
    x"1B",x"B7",x"C8",x"21",x"26",x"D6",x"CB",x"46", -- 0x0390
    x"36",x"00",x"28",x"02",x"EE",x"A0",x"C3",x"D6", -- 0x0398
    x"D5",x"3A",x"08",x"D6",x"2F",x"6F",x"AF",x"67", -- 0x03A0
    x"CB",x"7D",x"C0",x"7D",x"FE",x"0F",x"38",x"09", -- 0x03A8
    x"7D",x"D6",x"0B",x"6F",x"FE",x"0F",x"3E",x"20", -- 0x03B0
    x"D8",x"7D",x"FE",x"23",x"38",x"06",x"11",x"8E", -- 0x03B8
    x"1C",x"19",x"7E",x"C9",x"FE",x"13",x"20",x"0A", -- 0x03C0
    x"3A",x"24",x"D6",x"07",x"3E",x"0D",x"D0",x"3E", -- 0x03C8
    x"1B",x"C9",x"54",x"5D",x"29",x"19",x"11",x"5A", -- 0x03D0
    x"1C",x"19",x"46",x"EB",x"21",x"1E",x"D6",x"CB", -- 0x03D8
    x"7E",x"20",x"28",x"13",x"23",x"23",x"CB",x"7E", -- 0x03E0
    x"20",x"25",x"13",x"23",x"23",x"CB",x"7E",x"20", -- 0x03E8
    x"1E",x"78",x"2A",x"24",x"D6",x"FE",x"5C",x"38", -- 0x03F0
    x"08",x"C6",x"24",x"CB",x"7D",x"C8",x"C6",x"04", -- 0x03F8
    x"C9",x"CD",x"D0",x"D5",x"7C",x"AD",x"78",x"F8", -- 0x0400
    x"EE",x"20",x"C9",x"78",x"D6",x"40",x"C9",x"1A", -- 0x0408
    x"C9",x"4F",x"11",x"1E",x"D6",x"21",x"40",x"1C", -- 0x0410
    x"06",x"04",x"79",x"E6",x"3F",x"BE",x"23",x"20", -- 0x0418
    x"11",x"79",x"2F",x"12",x"07",x"30",x"16",x"EB", -- 0x0420
    x"23",x"3A",x"1E",x"D6",x"AE",x"77",x"AF",x"C3", -- 0x0428
    x"D9",x"D5",x"13",x"13",x"10",x"E4",x"EB",x"79", -- 0x0430
    x"FE",x"57",x"20",x"01",x"34",x"C3",x"5E",x"1B", -- 0x0438
    x"28",x"16",x"0F",x"19",x"E5",x"D5",x"CD",x"4C", -- 0x0440
    x"1C",x"D1",x"E1",x"C9",x"21",x"09",x"D6",x"7E", -- 0x0448
    x"B7",x"C8",x"E5",x"23",x"23",x"CD",x"51",x"1B", -- 0x0450
    x"7E",x"E1",x"35",x"B7",x"C9",x"52",x"34",x"24", -- 0x0458
    x"45",x"33",x"23",x"57",x"32",x"22",x"54",x"35", -- 0x0460
    x"25",x"51",x"31",x"21",x"46",x"7C",x"5E",x"44", -- 0x0468
    x"60",x"3D",x"53",x"2B",x"2B",x"47",x"5F",x"5F", -- 0x0470
    x"41",x"7E",x"2D",x"43",x"7F",x"3A",x"58",x"5C", -- 0x0478
    x"2F",x"5A",x"2A",x"2A",x"56",x"3B",x"3B",x"4A", -- 0x0480
    x"3E",x"3E",x"4B",x"7B",x"5B",x"4C",x"7D",x"5D", -- 0x0488
    x"48",x"3C",x"3C",x"FF",x"FF",x"FF",x"55",x"37", -- 0x0490
    x"27",x"49",x"38",x"28",x"4F",x"39",x"29",x"59", -- 0x0498
    x"36",x"26",x"50",x"30",x"40",x"4E",x"2C",x"2C", -- 0x04A0
    x"4D",x"2E",x"2E",x"5C",x"8C",x"88",x"42",x"3F", -- 0x04A8
    x"3F",x"82",x"81",x"80",x"83",x"20",x"FF",x"5D", -- 0x04B0
    x"8D",x"89",x"5F",x"8F",x"8B",x"FF",x"FF",x"FF", -- 0x04B8
    x"5E",x"8E",x"8A",x"1F",x"16",x"0F",x"1F",x"1F", -- 0x04C0
    x"00",x"01",x"0F",x"1F",x"1F",x"E5",x"D5",x"C5", -- 0x04C8
    x"F5",x"4F",x"21",x"2E",x"D6",x"E5",x"CB",x"D6", -- 0x04D0
    x"CB",x"46",x"C5",x"C4",x"C2",x"18",x"C1",x"CD", -- 0x04D8
    x"EA",x"1C",x"E1",x"CB",x"96",x"F1",x"C1",x"D1", -- 0x04E0
    x"E1",x"C9",x"2A",x"E3",x"D4",x"E5",x"21",x"F6", -- 0x04E8
    x"1C",x"22",x"E3",x"D4",x"79",x"C9",x"FE",x"20", -- 0x04F0
    x"30",x"1C",x"2A",x"C4",x"D4",x"87",x"5F",x"16", -- 0x04F8
    x"00",x"19",x"5E",x"23",x"56",x"D5",x"ED",x"5B", -- 0x0500
    x"34",x"D6",x"2A",x"36",x"D6",x"C9",x"26",x"00", -- 0x0508
    x"CD",x"BE",x"1E",x"6F",x"18",x"1D",x"F5",x"CD", -- 0x0510
    x"06",x"1D",x"3A",x"3A",x"D6",x"B7",x"C4",x"4D", -- 0x0518
    x"1D",x"2A",x"36",x"D6",x"F1",x"CD",x"37",x"1D", -- 0x0520
    x"CD",x"06",x"1D",x"2C",x"7D",x"BB",x"38",x"03", -- 0x0528
    x"32",x"3A",x"D6",x"22",x"36",x"D6",x"C9",x"47", -- 0x0530
    x"ED",x"5B",x"38",x"D6",x"19",x"E5",x"CD",x"4F", -- 0x0538
    x"1F",x"70",x"E1",x"78",x"C3",x"A6",x"D4",x"3A", -- 0x0540
    x"31",x"D6",x"B7",x"20",x"C3",x"CD",x"BE",x"1E", -- 0x0548
    x"6F",x"24",x"7C",x"BA",x"38",x"DD",x"25",x"22", -- 0x0550
    x"36",x"D6",x"21",x"00",x"00",x"4D",x"44",x"24", -- 0x0558
    x"15",x"28",x"2B",x"CD",x"68",x"1D",x"18",x"F5", -- 0x0560
    x"E5",x"D5",x"C5",x"E5",x"2A",x"38",x"D6",x"E5", -- 0x0568
    x"09",x"4B",x"D1",x"E3",x"19",x"D1",x"06",x"00", -- 0x0570
    x"E5",x"D5",x"C5",x"CD",x"4F",x"1F",x"EB",x"CD", -- 0x0578
    x"4F",x"1F",x"EB",x"ED",x"B0",x"C1",x"D1",x"E1", -- 0x0580
    x"CD",x"A9",x"D4",x"C3",x"E6",x"1C",x"CD",x"06", -- 0x0588
    x"1D",x"2E",x"00",x"7B",x"95",x"5F",x"C8",x"44", -- 0x0590
    x"4D",x"2A",x"38",x"D6",x"09",x"E5",x"43",x"CD", -- 0x0598
    x"4F",x"1F",x"AF",x"77",x"23",x"10",x"FC",x"E1", -- 0x05A0
    x"C3",x"AC",x"D4",x"24",x"7C",x"BA",x"D0",x"18", -- 0x05A8
    x"82",x"E5",x"D5",x"CD",x"93",x"1D",x"D1",x"E1", -- 0x05B0
    x"2E",x"00",x"24",x"7C",x"BA",x"38",x"F2",x"C9", -- 0x05B8
    x"CD",x"C8",x"1D",x"3E",x"20",x"CD",x"16",x"1D", -- 0x05C0
    x"CD",x"BE",x"1E",x"7C",x"B5",x"C8",x"CD",x"E2", -- 0x05C8
    x"1D",x"EF",x"C8",x"37",x"18",x"D9",x"CD",x"BE", -- 0x05D0
    x"1E",x"EF",x"C8",x"CD",x"09",x"1E",x"7C",x"BA", -- 0x05D8
    x"38",x"CD",x"7C",x"B5",x"C8",x"2D",x"F0",x"6B", -- 0x05E0
    x"2D",x"25",x"C9",x"E5",x"44",x"4D",x"CD",x"D6", -- 0x05E8
    x"1D",x"30",x"0C",x"EF",x"28",x"09",x"D5",x"1E", -- 0x05F0
    x"01",x"CD",x"68",x"1D",x"D1",x"18",x"ED",x"60", -- 0x05F8
    x"69",x"1E",x"01",x"CD",x"97",x"1D",x"E1",x"18", -- 0x0600
    x"A6",x"2C",x"7D",x"BB",x"D8",x"2E",x"00",x"24", -- 0x0608
    x"C9",x"CD",x"C8",x"1D",x"38",x"FB",x"C9",x"CD", -- 0x0610
    x"D6",x"1D",x"38",x"FB",x"C9",x"3E",x"09",x"CD", -- 0x0618
    x"16",x"1D",x"2A",x"36",x"D6",x"7D",x"E6",x"07", -- 0x0620
    x"3E",x"19",x"20",x"F3",x"C9",x"21",x"2E",x"D6", -- 0x0628
    x"CB",x"CE",x"C9",x"21",x"2E",x"D6",x"CB",x"8E", -- 0x0630
    x"C9",x"3E",x"AF",x"32",x"32",x"D6",x"C9",x"CF", -- 0x0638
    x"2A",x"34",x"D6",x"BC",x"D0",x"32",x"37",x"D6", -- 0x0640
    x"18",x"09",x"CF",x"2A",x"34",x"D6",x"BD",x"D0", -- 0x0648
    x"32",x"36",x"D6",x"18",x"69",x"CF",x"4F",x"3A", -- 0x0650
    x"29",x"D6",x"B9",x"C8",x"CD",x"B2",x"D4",x"EB", -- 0x0658
    x"21",x"31",x"D6",x"CD",x"70",x"1E",x"79",x"32", -- 0x0660
    x"29",x"D6",x"CD",x"B2",x"D4",x"11",x"31",x"D6", -- 0x0668
    x"C5",x"01",x"0A",x"00",x"ED",x"B0",x"C1",x"C9", -- 0x0670
    x"21",x"3B",x"D6",x"FE",x"08",x"D0",x"11",x"0A", -- 0x0678
    x"00",x"3D",x"F8",x"19",x"18",x"FB",x"CF",x"32", -- 0x0680
    x"2A",x"D6",x"CF",x"32",x"2B",x"D6",x"CF",x"32", -- 0x0688
    x"2C",x"D6",x"CF",x"32",x"2D",x"D6",x"2A",x"2A", -- 0x0690
    x"D6",x"EB",x"2A",x"2C",x"D6",x"ED",x"4B",x"E1", -- 0x0698
    x"D4",x"7C",x"B7",x"C8",x"82",x"3D",x"B8",x"D0", -- 0x06A0
    x"7D",x"B7",x"C8",x"83",x"3D",x"B9",x"D0",x"2A", -- 0x06A8
    x"2A",x"D6",x"22",x"38",x"D6",x"CD",x"0E",x"1D", -- 0x06B0
    x"2A",x"2C",x"D6",x"22",x"34",x"D6",x"AF",x"32", -- 0x06B8
    x"3A",x"D6",x"C9",x"21",x"FF",x"19",x"11",x"E0", -- 0x06C0
    x"D4",x"01",x"05",x"00",x"ED",x"B0",x"3E",x"FC", -- 0x06C8
    x"CD",x"FD",x"1E",x"3E",x"07",x"DF",x"11",x"D7", -- 0x06D0
    x"DF",x"12",x"DF",x"00",x"DF",x"00",x"DF",x"28", -- 0x06D8
    x"DF",x"15",x"3D",x"F2",x"D5",x"1E",x"C9",x"CF", -- 0x06E0
    x"FE",x"49",x"28",x"D7",x"21",x"27",x"D6",x"FE", -- 0x06E8
    x"53",x"28",x"14",x"FE",x"46",x"28",x"0D",x"FE", -- 0x06F0
    x"4C",x"C2",x"AF",x"D5",x"CF",x"0F",x"4F",x"06", -- 0x06F8
    x"40",x"ED",x"78",x"C9",x"CB",x"86",x"C9",x"CB", -- 0x0700
    x"C6",x"C9",x"44",x"4D",x"CD",x"17",x"1E",x"7C", -- 0x0708
    x"B8",x"20",x"0A",x"CD",x"33",x"1D",x"79",x"BD", -- 0x0710
    x"3E",x"20",x"D2",x"37",x"1D",x"C5",x"44",x"4D", -- 0x0718
    x"CD",x"E2",x"1D",x"D5",x"1E",x"01",x"CD",x"68", -- 0x0720
    x"1D",x"D1",x"C1",x"18",x"E2",x"EB",x"25",x"5D", -- 0x0728
    x"2E",x"00",x"7A",x"BC",x"D2",x"93",x"1D",x"44", -- 0x0730
    x"4D",x"25",x"CD",x"68",x"1D",x"18",x"F3",x"2E", -- 0x0738
    x"00",x"44",x"4D",x"7C",x"3C",x"BA",x"D2",x"93", -- 0x0740
    x"1D",x"24",x"CD",x"68",x"1D",x"18",x"F2",x"D5", -- 0x0748
    x"E5",x"6C",x"26",x"00",x"CD",x"A3",x"D4",x"D1", -- 0x0750
    x"16",x"00",x"19",x"ED",x"5B",x"BC",x"D4",x"19", -- 0x0758
    x"D1",x"C9",x"29",x"29",x"29",x"54",x"5D",x"29", -- 0x0760
    x"29",x"19",x"C9",x"A3",x"D5",x"3F",x"1E",x"4A", -- 0x0768
    x"1E",x"39",x"1E",x"3A",x"1E",x"11",x"1E",x"17", -- 0x0770
    x"1E",x"AD",x"19",x"C0",x"1D",x"1D",x"1E",x"51", -- 0x0778
    x"1D",x"A6",x"D5",x"A9",x"D5",x"4D",x"1D",x"2D", -- 0x0780
    x"1E",x"33",x"1E",x"AC",x"D5",x"55",x"1E",x"86", -- 0x0788
    x"1E",x"EB",x"1D",x"0A",x"1F",x"3F",x"1F",x"2D", -- 0x0790
    x"1F",x"13",x"18",x"C8",x"1D",x"D6",x"1D",x"AB", -- 0x0798
    x"1D",x"E7",x"1E",x"0E",x"1D",x"10",x"1D",x"93", -- 0x07A0
    x"1D",x"B1",x"1D",x"E5",x"D5",x"C5",x"21",x"8B", -- 0x07A8
    x"D6",x"06",x"0C",x"36",x"00",x"23",x"10",x"FB", -- 0x07B0
    x"FE",x"80",x"30",x"22",x"D6",x"21",x"D4",x"A6", -- 0x07B8
    x"20",x"C1",x"D1",x"E1",x"F7",x"11",x"8B",x"D6", -- 0x07C0
    x"01",x"00",x"0C",x"3A",x"32",x"D6",x"B7",x"28", -- 0x07C8
    x"01",x"0D",x"1A",x"13",x"A9",x"77",x"CB",x"05", -- 0x07D0
    x"2C",x"CB",x"0D",x"10",x"F5",x"C9",x"FE",x"C0", -- 0x07D8
    x"30",x"23",x"D6",x"80",x"5F",x"16",x"00",x"2A", -- 0x07E0
    x"00",x"D6",x"7D",x"B4",x"28",x"D3",x"EB",x"29", -- 0x07E8
    x"29",x"44",x"4D",x"29",x"09",x"19",x"11",x"8B", -- 0x07F0
    x"D6",x"06",x"0C",x"CD",x"12",x"D5",x"23",x"12", -- 0x07F8
    x"13",x"10",x"F8",x"18",x"BC",x"0E",x"3F",x"FE", -- 0x0800
    x"E0",x"38",x"02",x"0E",x"1F",x"E6",x"1F",x"5F", -- 0x0808
    x"16",x"00",x"21",x"CD",x"27",x"19",x"7E",x"B7", -- 0x0810
    x"28",x"A7",x"F5",x"E6",x"1F",x"28",x"04",x"81", -- 0x0818
    x"CD",x"A6",x"20",x"F1",x"0F",x"0F",x"0F",x"0F", -- 0x0820
    x"E6",x"0E",x"5F",x"16",x"00",x"21",x"BD",x"27", -- 0x0828
    x"19",x"11",x"94",x"D6",x"01",x"02",x"00",x"ED", -- 0x0830
    x"B0",x"18",x"86",x"F7",x"06",x"0C",x"7E",x"2F", -- 0x0838
    x"77",x"CB",x"05",x"2C",x"CB",x"0D",x"10",x"F6", -- 0x0840
    x"21",x"2E",x"D6",x"7E",x"EE",x"01",x"77",x"C9", -- 0x0848
    x"E5",x"D5",x"C5",x"21",x"8B",x"D6",x"11",x"8C", -- 0x0850
    x"D6",x"01",x"0B",x"00",x"3A",x"32",x"D6",x"B7", -- 0x0858
    x"28",x"02",x"3E",x"FF",x"77",x"ED",x"B0",x"C1", -- 0x0860
    x"D1",x"E1",x"F7",x"EB",x"E5",x"D5",x"21",x"8B", -- 0x0868
    x"D6",x"01",x"06",x"00",x"ED",x"B0",x"7B",x"D6", -- 0x0870
    x"85",x"5F",x"0E",x"06",x"ED",x"B0",x"D1",x"E1", -- 0x0878
    x"15",x"2D",x"20",x"E8",x"C9",x"F7",x"EB",x"F7", -- 0x0880
    x"EB",x"41",x"E5",x"D5",x"C5",x"01",x"06",x"00", -- 0x0888
    x"ED",x"B0",x"7D",x"D6",x"85",x"6F",x"7B",x"D6", -- 0x0890
    x"85",x"5F",x"0E",x"06",x"ED",x"B0",x"C1",x"D1", -- 0x0898
    x"E1",x"25",x"15",x"10",x"E5",x"C9",x"5F",x"16", -- 0x08A0
    x"00",x"62",x"6B",x"29",x"19",x"29",x"19",x"11", -- 0x08A8
    x"24",x"25",x"19",x"11",x"8D",x"D6",x"01",x"07", -- 0x08B0
    x"00",x"CB",x"46",x"28",x"02",x"1B",x"1B",x"D5", -- 0x08B8
    x"ED",x"B0",x"FE",x"49",x"20",x"04",x"13",x"3E", -- 0x08C0
    x"18",x"12",x"E1",x"CB",x"86",x"C9",x"CD",x"C1", -- 0x08C8
    x"D5",x"CD",x"12",x"D5",x"FE",x"23",x"20",x"03", -- 0x08D0
    x"CB",x"D0",x"23",x"CB",x"E8",x"C5",x"D5",x"11", -- 0x08D8
    x"97",x"D6",x"01",x"20",x"0C",x"CD",x"0A",x"21", -- 0x08E0
    x"23",x"28",x"01",x"E3",x"06",x"03",x"3E",x"2E", -- 0x08E8
    x"12",x"13",x"CD",x"0A",x"21",x"EB",x"D1",x"71", -- 0x08F0
    x"23",x"71",x"23",x"36",x"31",x"23",x"AF",x"77", -- 0x08F8
    x"23",x"77",x"23",x"77",x"23",x"C1",x"71",x"23", -- 0x0900
    x"70",x"C9",x"CD",x"12",x"D5",x"23",x"FE",x"2E", -- 0x0908
    x"F5",x"28",x"03",x"B9",x"30",x"02",x"2B",x"79", -- 0x0910
    x"12",x"13",x"F1",x"10",x"ED",x"C9",x"CD",x"AD", -- 0x0918
    x"22",x"21",x"97",x"D6",x"AF",x"CD",x"C9",x"22", -- 0x0920
    x"CD",x"E2",x"22",x"21",x"AF",x"D6",x"E5",x"01", -- 0x0928
    x"17",x"00",x"3E",x"48",x"CD",x"EA",x"22",x"E1", -- 0x0930
    x"20",x"58",x"11",x"97",x"D6",x"06",x"13",x"1A", -- 0x0938
    x"FE",x"20",x"20",x"06",x"80",x"FE",x"24",x"30", -- 0x0940
    x"04",x"90",x"BE",x"20",x"39",x"23",x"13",x"10", -- 0x0948
    x"EE",x"2A",x"BE",x"D4",x"ED",x"4B",x"C3",x"D6", -- 0x0950
    x"3E",x"44",x"CD",x"EA",x"22",x"20",x"33",x"21", -- 0x0958
    x"AF",x"D6",x"11",x"97",x"D6",x"01",x"10",x"00", -- 0x0960
    x"ED",x"B0",x"DF",x"1D",x"DF",x"1E",x"21",x"AE", -- 0x0968
    x"D6",x"CB",x"DE",x"CB",x"46",x"C4",x"D6",x"22", -- 0x0970
    x"CD",x"B8",x"22",x"F1",x"C1",x"D1",x"E1",x"D9", -- 0x0978
    x"08",x"AF",x"C1",x"D1",x"E1",x"C9",x"21",x"AF", -- 0x0980
    x"D6",x"3E",x"14",x"CD",x"C9",x"22",x"DF",x"07", -- 0x0988
    x"18",x"96",x"21",x"CE",x"23",x"06",x"0F",x"3E", -- 0x0990
    x"14",x"CD",x"CB",x"22",x"18",x"F0",x"CD",x"C4", -- 0x0998
    x"D5",x"E5",x"21",x"AE",x"D6",x"CB",x"56",x"20", -- 0x09A0
    x"35",x"CB",x"5E",x"28",x"24",x"2A",x"C3",x"D6", -- 0x09A8
    x"7C",x"B5",x"28",x"17",x"2B",x"22",x"C3",x"D6", -- 0x09B0
    x"2A",x"AB",x"D6",x"23",x"22",x"AB",x"D6",x"2B", -- 0x09B8
    x"D5",x"ED",x"5B",x"BE",x"D4",x"19",x"D1",x"AF", -- 0x09C0
    x"7E",x"E1",x"C9",x"3A",x"C2",x"D6",x"B7",x"3E", -- 0x09C8
    x"00",x"CC",x"1E",x"21",x"21",x"00",x"00",x"22", -- 0x09D0
    x"AB",x"D6",x"28",x"D1",x"E1",x"C9",x"F3",x"C5", -- 0x09D8
    x"3E",x"04",x"D3",x"03",x"26",x"FF",x"CB",x"76", -- 0x09E0
    x"28",x"FC",x"CB",x"76",x"20",x"FC",x"0E",x"80", -- 0x09E8
    x"3A",x"C6",x"D4",x"47",x"10",x"FE",x"3A",x"C7", -- 0x09F0
    x"D4",x"47",x"7E",x"07",x"07",x"CB",x"19",x"30", -- 0x09F8
    x"F3",x"10",x"FE",x"7E",x"2F",x"CB",x"77",x"3A", -- 0x0A00
    x"27",x"D6",x"D3",x"03",x"79",x"C1",x"E1",x"C9", -- 0x0A08
    x"6F",x"26",x"FF",x"F3",x"C5",x"D5",x"4D",x"ED", -- 0x0A10
    x"5B",x"C8",x"D4",x"AF",x"D3",x"03",x"9F",x"E6", -- 0x0A18
    x"06",x"F6",x"09",x"D3",x"0A",x"43",x"10",x"FE", -- 0x0A20
    x"CB",x"2C",x"CB",x"1D",x"15",x"20",x"EF",x"D1", -- 0x0A28
    x"18",x"D5",x"CD",x"C7",x"D5",x"E5",x"21",x"AE", -- 0x0A30
    x"D6",x"CB",x"E6",x"CB",x"56",x"20",x"D1",x"2A", -- 0x0A38
    x"AB",x"D6",x"CB",x"54",x"20",x"0F",x"23",x"22", -- 0x0A40
    x"AB",x"D6",x"2B",x"D5",x"ED",x"5B",x"BE",x"D4", -- 0x0A48
    x"19",x"D1",x"77",x"E1",x"C9",x"F5",x"CD",x"74", -- 0x0A50
    x"22",x"F1",x"18",x"E3",x"CD",x"CA",x"D5",x"E5", -- 0x0A58
    x"21",x"AE",x"D6",x"CB",x"66",x"28",x"A7",x"CB", -- 0x0A60
    x"56",x"21",x"00",x"FE",x"20",x"A5",x"E1",x"3E", -- 0x0A68
    x"FF",x"32",x"AA",x"D6",x"CD",x"AD",x"22",x"CD", -- 0x0A70
    x"E2",x"22",x"F3",x"21",x"AE",x"D6",x"01",x"80", -- 0x0A78
    x"00",x"7E",x"E6",x"22",x"CB",x"AE",x"28",x"01", -- 0x0A80
    x"04",x"CD",x"82",x"23",x"21",x"97",x"D6",x"01", -- 0x0A88
    x"17",x"00",x"3E",x"48",x"CD",x"6A",x"23",x"2A", -- 0x0A90
    x"BE",x"D4",x"ED",x"4B",x"AB",x"D6",x"3E",x"44", -- 0x0A98
    x"CD",x"6A",x"23",x"FB",x"21",x"00",x"00",x"22", -- 0x0AA0
    x"AB",x"D6",x"C3",x"6E",x"21",x"E3",x"D5",x"C5", -- 0x0AA8
    x"D9",x"08",x"E5",x"D5",x"C5",x"F5",x"D9",x"E9", -- 0x0AB0
    x"21",x"A9",x"D6",x"34",x"7E",x"FE",x"31",x"38", -- 0x0AB8
    x"FA",x"FE",x"3A",x"D8",x"36",x"30",x"2B",x"18", -- 0x0AC0
    x"F2",x"06",x"13",x"DF",x"02",x"D7",x"7E",x"23", -- 0x0AC8
    x"D7",x"10",x"FB",x"DF",x"1E",x"C9",x"3A",x"28", -- 0x0AD0
    x"D6",x"E6",x"EE",x"3C",x"32",x"28",x"D6",x"D3", -- 0x0AD8
    x"0A",x"C9",x"3A",x"28",x"D6",x"F6",x"11",x"3D", -- 0x0AE0
    x"18",x"F2",x"32",x"C6",x"D6",x"3A",x"27",x"D6", -- 0x0AE8
    x"F5",x"C5",x"E5",x"37",x"08",x"21",x"27",x"D6", -- 0x0AF0
    x"7E",x"F6",x"05",x"77",x"D3",x"03",x"11",x"32", -- 0x0AF8
    x"00",x"26",x"FF",x"FB",x"76",x"F3",x"3D",x"D3", -- 0x0B00
    x"03",x"1B",x"CD",x"52",x"23",x"38",x"FA",x"CB", -- 0x0B08
    x"7A",x"28",x"E0",x"57",x"08",x"D9",x"CD",x"3A", -- 0x0B10
    x"23",x"2A",x"C6",x"D6",x"BD",x"20",x"D4",x"08", -- 0x0B18
    x"16",x"00",x"E1",x"C1",x"CD",x"3A",x"23",x"77", -- 0x0B20
    x"82",x"57",x"ED",x"A1",x"EA",x"24",x"23",x"CD", -- 0x0B28
    x"3A",x"23",x"BA",x"21",x"27",x"D6",x"C1",x"70", -- 0x0B30
    x"FF",x"C9",x"D9",x"CD",x"52",x"23",x"DC",x"52", -- 0x0B38
    x"23",x"1E",x"80",x"CD",x"52",x"23",x"DC",x"52", -- 0x0B40
    x"23",x"AA",x"07",x"CB",x"1B",x"30",x"F4",x"7B", -- 0x0B48
    x"D9",x"C9",x"06",x"0E",x"CD",x"C2",x"23",x"06", -- 0x0B50
    x"25",x"7E",x"AD",x"FA",x"B9",x"23",x"10",x"F9", -- 0x0B58
    x"D1",x"08",x"38",x"8F",x"D1",x"20",x"8C",x"B4", -- 0x0B60
    x"18",x"C9",x"08",x"D9",x"11",x"00",x"03",x"37", -- 0x0B68
    x"CD",x"A5",x"23",x"1B",x"7A",x"B3",x"20",x"F7", -- 0x0B70
    x"CD",x"A5",x"23",x"08",x"D9",x"CD",x"92",x"23", -- 0x0B78
    x"16",x"00",x"7E",x"CD",x"92",x"23",x"7E",x"82", -- 0x0B80
    x"57",x"ED",x"A1",x"EA",x"82",x"23",x"7A",x"CD", -- 0x0B88
    x"92",x"23",x"D9",x"5F",x"1F",x"3F",x"CD",x"A5", -- 0x0B90
    x"23",x"37",x"CB",x"1B",x"CD",x"A5",x"23",x"CB", -- 0x0B98
    x"3B",x"20",x"F9",x"D9",x"C9",x"9F",x"E6",x"08", -- 0x0BA0
    x"6F",x"06",x"19",x"CD",x"C2",x"23",x"7D",x"D3", -- 0x0BA8
    x"03",x"EE",x"08",x"06",x"1F",x"10",x"FE",x"D3", -- 0x0BB0
    x"03",x"3E",x"1A",x"B8",x"ED",x"5F",x"4F",x"7E", -- 0x0BB8
    x"6F",x"C9",x"ED",x"5F",x"91",x"E6",x"7F",x"CB", -- 0x0BC0
    x"3F",x"90",x"3C",x"20",x"FD",x"C9",x"43",x"68", -- 0x0BC8
    x"79",x"62",x"61",x"20",x"70",x"D2",x"69",x"20", -- 0x0BD0
    x"C3",x"74",x"65",x"6E",x"C9",x"E5",x"01",x"DE", -- 0x0BD8
    x"23",x"C5",x"CD",x"1E",x"24",x"FE",x"80",x"28", -- 0x0BE0
    x"16",x"FE",x"83",x"28",x"16",x"FE",x"0D",x"28", -- 0x0BE8
    x"17",x"FE",x"84",x"28",x"07",x"FE",x"1F",x"C2", -- 0x0BF0
    x"B8",x"D5",x"D7",x"C9",x"DF",x"1C",x"C9",x"DF", -- 0x0BF8
    x"17",x"18",x"02",x"DF",x"0A",x"C3",x"A5",x"24", -- 0x0C00
    x"C1",x"C1",x"C5",x"2A",x"C8",x"D6",x"EF",x"02", -- 0x0C08
    x"28",x"06",x"03",x"CD",x"09",x"1E",x"18",x"F6", -- 0x0C10
    x"DF",x"06",x"DF",x"0D",x"E1",x"C9",x"DF",x"0E", -- 0x0C18
    x"2A",x"36",x"D6",x"E5",x"DF",x"05",x"2A",x"36", -- 0x0C20
    x"D6",x"22",x"C8",x"D6",x"DF",x"06",x"2A",x"36", -- 0x0C28
    x"D6",x"22",x"CA",x"D6",x"E1",x"E7",x"01",x"36", -- 0x0C30
    x"24",x"C5",x"CD",x"06",x"1D",x"CD",x"AC",x"1A", -- 0x0C38
    x"4F",x"E6",x"7F",x"FE",x"20",x"79",x"DA",x"C6", -- 0x0C40
    x"24",x"3A",x"CA",x"D6",x"3C",x"BB",x"38",x"2B", -- 0x0C48
    x"3A",x"CB",x"D6",x"3C",x"BA",x"38",x"16",x"3A", -- 0x0C50
    x"C9",x"D6",x"B7",x"C8",x"E5",x"DF",x"01",x"AF", -- 0x0C58
    x"D7",x"DF",x"15",x"21",x"C9",x"D6",x"35",x"21", -- 0x0C60
    x"CB",x"D6",x"35",x"E1",x"25",x"E5",x"2A",x"CA", -- 0x0C68
    x"D6",x"CD",x"09",x"1E",x"EF",x"28",x"03",x"E7", -- 0x0C70
    x"DF",x"16",x"E1",x"E5",x"2A",x"CA",x"D6",x"CD", -- 0x0C78
    x"09",x"1E",x"22",x"CA",x"D6",x"E1",x"E7",x"DF", -- 0x0C80
    x"14",x"79",x"D7",x"7D",x"3C",x"BB",x"D8",x"DF", -- 0x0C88
    x"0D",x"C9",x"3A",x"C9",x"D6",x"BC",x"28",x"52", -- 0x0C90
    x"DF",x"17",x"C9",x"3A",x"CB",x"D6",x"94",x"28", -- 0x0C98
    x"49",x"DF",x"1A",x"3D",x"C0",x"2A",x"36",x"D6", -- 0x0CA0
    x"EF",x"C0",x"E7",x"7D",x"B7",x"C8",x"CD",x"E2", -- 0x0CA8
    x"1D",x"18",x"F5",x"E5",x"E7",x"DF",x"1E",x"2E", -- 0x0CB0
    x"00",x"3A",x"CB",x"D6",x"24",x"BC",x"30",x"F4", -- 0x0CB8
    x"E1",x"22",x"CA",x"D6",x"E7",x"C9",x"FE",x"81", -- 0x0CC0
    x"28",x"23",x"FE",x"82",x"28",x"2A",x"FE",x"1C", -- 0x0CC8
    x"28",x"3C",x"FE",x"1D",x"28",x"2F",x"FE",x"85", -- 0x0CD0
    x"28",x"44",x"FE",x"86",x"28",x"43",x"FE",x"1E", -- 0x0CD8
    x"28",x"D1",x"FE",x"80",x"28",x"AC",x"FE",x"83", -- 0x0CE0
    x"28",x"B1",x"79",x"C1",x"C9",x"DF",x"18",x"C9", -- 0x0CE8
    x"7D",x"B7",x"C0",x"3A",x"C9",x"D6",x"BC",x"C9", -- 0x0CF0
    x"DF",x"19",x"C9",x"3A",x"CB",x"D6",x"BC",x"C0", -- 0x0CF8
    x"3A",x"CA",x"D6",x"BD",x"C9",x"CD",x"F0",x"24", -- 0x0D00
    x"C8",x"DF",x"18",x"2A",x"36",x"D6",x"CD",x"FB", -- 0x0D08
    x"24",x"C8",x"DF",x"13",x"2A",x"CA",x"D6",x"CD", -- 0x0D10
    x"E2",x"1D",x"22",x"CA",x"D6",x"C9",x"DF",x"05", -- 0x0D18
    x"C9",x"DF",x"06",x"C9",x"30",x"00",x"30",x"30", -- 0x0D20
    x"78",x"78",x"30",x"00",x"00",x"00",x"00",x"6C", -- 0x0D28
    x"6C",x"6C",x"6C",x"6C",x"FE",x"6C",x"FE",x"6C", -- 0x0D30
    x"6C",x"30",x"F8",x"0C",x"78",x"C0",x"7C",x"30", -- 0x0D38
    x"C6",x"66",x"30",x"18",x"CC",x"C6",x"00",x"76", -- 0x0D40
    x"CC",x"DC",x"76",x"38",x"6C",x"38",x"00",x"00", -- 0x0D48
    x"00",x"00",x"60",x"30",x"30",x"18",x"30",x"60", -- 0x0D50
    x"60",x"60",x"30",x"18",x"60",x"30",x"18",x"18", -- 0x0D58
    x"18",x"30",x"60",x"00",x"6C",x"38",x"FE",x"38", -- 0x0D60
    x"6C",x"00",x"00",x"30",x"30",x"FC",x"30",x"30", -- 0x0D68
    x"00",x"61",x"30",x"30",x"00",x"00",x"00",x"00", -- 0x0D70
    x"00",x"00",x"00",x"FC",x"00",x"00",x"00",x"30", -- 0x0D78
    x"30",x"00",x"00",x"00",x"00",x"00",x"00",x"C0", -- 0x0D80
    x"60",x"30",x"18",x"0C",x"06",x"78",x"CC",x"EC", -- 0x0D88
    x"FC",x"DC",x"CC",x"78",x"FC",x"30",x"30",x"30", -- 0x0D90
    x"F0",x"70",x"30",x"FC",x"CC",x"60",x"38",x"0C", -- 0x0D98
    x"CC",x"78",x"78",x"CC",x"0C",x"38",x"0C",x"CC", -- 0x0DA0
    x"78",x"1E",x"0C",x"FE",x"CC",x"6C",x"3C",x"1C", -- 0x0DA8
    x"78",x"CC",x"0C",x"0C",x"F8",x"C0",x"FC",x"78", -- 0x0DB0
    x"CC",x"CC",x"F8",x"C0",x"60",x"38",x"30",x"30", -- 0x0DB8
    x"30",x"7C",x"18",x"CC",x"FC",x"78",x"CC",x"CC", -- 0x0DC0
    x"78",x"CC",x"CC",x"78",x"70",x"18",x"0C",x"7C", -- 0x0DC8
    x"CC",x"CC",x"78",x"30",x"30",x"00",x"00",x"30", -- 0x0DD0
    x"30",x"00",x"61",x"30",x"30",x"00",x"00",x"30", -- 0x0DD8
    x"30",x"0C",x"18",x"30",x"60",x"30",x"18",x"0C", -- 0x0DE0
    x"00",x"FC",x"00",x"00",x"FC",x"00",x"00",x"60", -- 0x0DE8
    x"30",x"18",x"0C",x"18",x"30",x"60",x"30",x"00", -- 0x0DF0
    x"30",x"18",x"0C",x"CC",x"78",x"7E",x"C0",x"DE", -- 0x0DF8
    x"D6",x"D6",x"C6",x"7C",x"C6",x"C6",x"FE",x"C6", -- 0x0E00
    x"C6",x"6C",x"38",x"FC",x"66",x"66",x"7C",x"66", -- 0x0E08
    x"66",x"FC",x"7C",x"C6",x"C0",x"C0",x"C0",x"C6", -- 0x0E10
    x"7C",x"FC",x"66",x"66",x"66",x"66",x"66",x"FC", -- 0x0E18
    x"FE",x"62",x"68",x"78",x"68",x"62",x"FE",x"F0", -- 0x0E20
    x"60",x"68",x"78",x"68",x"62",x"FE",x"7C",x"C6", -- 0x0E28
    x"CE",x"C0",x"C0",x"C6",x"7C",x"C6",x"C6",x"C6", -- 0x0E30
    x"FE",x"C6",x"C6",x"C6",x"3C",x"18",x"18",x"18", -- 0x0E38
    x"18",x"18",x"3C",x"78",x"CC",x"CC",x"0C",x"0C", -- 0x0E40
    x"0C",x"1E",x"E6",x"66",x"6C",x"78",x"6C",x"66", -- 0x0E48
    x"E6",x"FE",x"66",x"60",x"60",x"60",x"60",x"F0", -- 0x0E50
    x"C6",x"C6",x"D6",x"FE",x"FE",x"EE",x"C6",x"C6", -- 0x0E58
    x"C6",x"CE",x"DE",x"F6",x"E6",x"C6",x"7C",x"C6", -- 0x0E60
    x"C6",x"C6",x"C6",x"C6",x"7C",x"F0",x"60",x"60", -- 0x0E68
    x"7C",x"66",x"66",x"FC",x"0E",x"7C",x"DE",x"C6", -- 0x0E70
    x"C6",x"C6",x"7C",x"E6",x"66",x"6C",x"7C",x"66", -- 0x0E78
    x"66",x"FC",x"7C",x"C6",x"06",x"7C",x"C0",x"C6", -- 0x0E80
    x"7C",x"78",x"30",x"30",x"30",x"30",x"B4",x"FC", -- 0x0E88
    x"7C",x"C6",x"C6",x"C6",x"C6",x"C6",x"C6",x"10", -- 0x0E90
    x"38",x"6C",x"C6",x"C6",x"C6",x"C6",x"C6",x"EE", -- 0x0E98
    x"FE",x"D6",x"C6",x"C6",x"C6",x"C6",x"6C",x"38", -- 0x0EA0
    x"38",x"6C",x"C6",x"C6",x"78",x"30",x"30",x"78", -- 0x0EA8
    x"CC",x"CC",x"CC",x"FE",x"66",x"32",x"18",x"8C", -- 0x0EB0
    x"C6",x"FE",x"78",x"60",x"60",x"60",x"60",x"60", -- 0x0EB8
    x"78",x"00",x"06",x"0C",x"18",x"30",x"60",x"C0", -- 0x0EC0
    x"78",x"18",x"18",x"18",x"18",x"18",x"78",x"30", -- 0x0EC8
    x"30",x"30",x"30",x"FC",x"78",x"30",x"FF",x"00", -- 0x0ED0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0ED8
    x"00",x"18",x"30",x"30",x"76",x"CC",x"7C",x"0C", -- 0x0EE0
    x"78",x"00",x"00",x"DC",x"66",x"66",x"66",x"7C", -- 0x0EE8
    x"60",x"E0",x"7C",x"C6",x"C0",x"C6",x"7C",x"00", -- 0x0EF0
    x"00",x"76",x"CC",x"CC",x"CC",x"7C",x"0C",x"1C", -- 0x0EF8
    x"7C",x"C0",x"FE",x"C6",x"7C",x"00",x"00",x"78", -- 0x0F00
    x"30",x"30",x"78",x"30",x"36",x"1C",x"F9",x"0C", -- 0x0F08
    x"7C",x"CC",x"CC",x"CC",x"76",x"E6",x"66",x"66", -- 0x0F10
    x"76",x"6C",x"60",x"E0",x"78",x"30",x"30",x"30", -- 0x0F18
    x"70",x"00",x"30",x"71",x"18",x"18",x"18",x"18", -- 0x0F20
    x"18",x"38",x"E6",x"6C",x"78",x"6C",x"66",x"60", -- 0x0F28
    x"E0",x"78",x"30",x"30",x"30",x"30",x"30",x"70", -- 0x0F30
    x"D6",x"D6",x"D6",x"FE",x"CC",x"00",x"00",x"C6", -- 0x0F38
    x"C6",x"C6",x"C6",x"FC",x"00",x"00",x"7C",x"C6", -- 0x0F40
    x"C6",x"C6",x"7C",x"00",x"00",x"F1",x"60",x"7C", -- 0x0F48
    x"66",x"66",x"66",x"DC",x"1F",x"0C",x"7C",x"CC", -- 0x0F50
    x"CC",x"CC",x"76",x"F0",x"60",x"66",x"76",x"DC", -- 0x0F58
    x"00",x"00",x"FC",x"06",x"7C",x"C0",x"7E",x"00", -- 0x0F60
    x"00",x"18",x"34",x"30",x"30",x"78",x"30",x"30", -- 0x0F68
    x"76",x"CC",x"CC",x"CC",x"CC",x"00",x"00",x"38", -- 0x0F70
    x"6C",x"C6",x"C6",x"C6",x"00",x"00",x"6C",x"FE", -- 0x0F78
    x"FE",x"D6",x"C6",x"00",x"00",x"C6",x"6C",x"38", -- 0x0F80
    x"6C",x"C6",x"00",x"00",x"7D",x"06",x"7E",x"C6", -- 0x0F88
    x"C6",x"C6",x"C6",x"FE",x"62",x"10",x"8C",x"FE", -- 0x0F90
    x"00",x"00",x"1C",x"30",x"30",x"E0",x"30",x"30", -- 0x0F98
    x"1C",x"18",x"18",x"18",x"00",x"18",x"18",x"18", -- 0x0FA0
    x"E0",x"30",x"30",x"1C",x"30",x"30",x"E0",x"00", -- 0x0FA8
    x"00",x"00",x"00",x"00",x"DC",x"76",x"AA",x"55", -- 0x0FB0
    x"AA",x"55",x"AA",x"55",x"AA",x"18",x"0C",x"18", -- 0x0FB8
    x"66",x"66",x"33",x"30",x"18",x"30",x"30",x"82", -- 0x0FC0
    x"7C",x"30",x"CC",x"60",x"C0",x"60",x"01",x"A2", -- 0x0FC8
    x"23",x"C4",x"C5",x"12",x"A8",x"55",x"09",x"95", -- 0x0FD0
    x"0C",x"2C",x"4F",x"CE",x"0F",x"AF",x"41",x"D2", -- 0x0FD8
    x"D3",x"D4",x"75",x"2F",x"65",x"E1",x"79",x"DA", -- 0x0FE0
    x"A7",x"C0",x"B0",x"80",x"B3",x"32",x"2E",x"37", -- 0x0FE8
    x"28",x"43",x"29",x"31",x"39",x"38",x"37",x"20", -- 0x0FF0
    x"56",x"69",x"4C",x"69",x"53",x"6F",x"66",x"74"  -- 0x0FF8
  );

begin

  p_rom : process
  begin
    wait until rising_edge(CLK);
    if (ENA = '1') then
       DATA <= ROM(to_integer(unsigned(ADDR)));
    end if;
  end process;
end RTL;
