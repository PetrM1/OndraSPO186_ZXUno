-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
--  
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity OndraSD_ZPU_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end OndraSD_ZPU_ROM;

architecture arch of OndraSD_ZPU_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
( 

0 => x"0b0b0b88", 
1 => x"e5040000", 
2 => x"00000000", 
3 => x"00000000", 
4 => x"00000000", 
5 => x"00000000", 
6 => x"00000000", 
7 => x"00000000", 
8 => x"88088c08", 
9 => x"90080b0b", 
10 => x"0b88e108", 
11 => x"2d900c8c", 
12 => x"0c880c04", 
13 => x"00000000", 
14 => x"00000000", 
15 => x"00000000", 
16 => x"71fd0608", 
17 => x"72830609", 
18 => x"81058205", 
19 => x"832b2a83", 
20 => x"ffff0652", 
21 => x"04000000", 
22 => x"00000000", 
23 => x"00000000", 
24 => x"71fd0608", 
25 => x"83ffff73", 
26 => x"83060981", 
27 => x"05820583", 
28 => x"2b2b0906", 
29 => x"7383ffff", 
30 => x"0b0b0b0b", 
31 => x"83a50400", 
32 => x"72098105", 
33 => x"72057373", 
34 => x"09060906", 
35 => x"73097306", 
36 => x"070a8106", 
37 => x"53510400", 
38 => x"00000000", 
39 => x"00000000", 
40 => x"72722473", 
41 => x"732e0753", 
42 => x"51040000", 
43 => x"00000000", 
44 => x"00000000", 
45 => x"00000000", 
46 => x"00000000", 
47 => x"00000000", 
48 => x"71737109", 
49 => x"71068106", 
50 => x"09810572", 
51 => x"0a100a72", 
52 => x"0a100a31", 
53 => x"050a8106", 
54 => x"51515351", 
55 => x"04000000", 
56 => x"72722673", 
57 => x"732e0753", 
58 => x"51040000", 
59 => x"00000000", 
60 => x"00000000", 
61 => x"00000000", 
62 => x"00000000", 
63 => x"00000000", 
64 => x"00000000", 
65 => x"00000000", 
66 => x"00000000", 
67 => x"00000000", 
68 => x"00000000", 
69 => x"00000000", 
70 => x"00000000", 
71 => x"00000000", 
72 => x"0b0b0b88", 
73 => x"ba040000", 
74 => x"00000000", 
75 => x"00000000", 
76 => x"00000000", 
77 => x"00000000", 
78 => x"00000000", 
79 => x"00000000", 
80 => x"720a722b", 
81 => x"0a535104", 
82 => x"00000000", 
83 => x"00000000", 
84 => x"00000000", 
85 => x"00000000", 
86 => x"00000000", 
87 => x"00000000", 
88 => x"72729f06", 
89 => x"0981050b", 
90 => x"0b0b889f", 
91 => x"05040000", 
92 => x"00000000", 
93 => x"00000000", 
94 => x"00000000", 
95 => x"00000000", 
96 => x"72722aff", 
97 => x"739f062a", 
98 => x"0974090a", 
99 => x"8106ff05", 
100 => x"06075351", 
101 => x"04000000", 
102 => x"00000000", 
103 => x"00000000", 
104 => x"71715351", 
105 => x"04067383", 
106 => x"06098105", 
107 => x"8205832b", 
108 => x"0b2b0772", 
109 => x"fc060c51", 
110 => x"51040000", 
111 => x"00000000", 
112 => x"72098105", 
113 => x"72050970", 
114 => x"81050906", 
115 => x"0a810653", 
116 => x"51040000", 
117 => x"00000000", 
118 => x"00000000", 
119 => x"00000000", 
120 => x"72098105", 
121 => x"72050970", 
122 => x"81050906", 
123 => x"0a098106", 
124 => x"53510400", 
125 => x"00000000", 
126 => x"00000000", 
127 => x"00000000", 
128 => x"71098105", 
129 => x"52040000", 
130 => x"00000000", 
131 => x"00000000", 
132 => x"00000000", 
133 => x"00000000", 
134 => x"00000000", 
135 => x"00000000", 
136 => x"72720981", 
137 => x"05055351", 
138 => x"04000000", 
139 => x"00000000", 
140 => x"00000000", 
141 => x"00000000", 
142 => x"00000000", 
143 => x"00000000", 
144 => x"72097206", 
145 => x"73730906", 
146 => x"07535104", 
147 => x"00000000", 
148 => x"00000000", 
149 => x"00000000", 
150 => x"00000000", 
151 => x"00000000", 
152 => x"71fc0608", 
153 => x"72830609", 
154 => x"81058305", 
155 => x"1010102a", 
156 => x"81ff0652", 
157 => x"04000000", 
158 => x"00000000", 
159 => x"00000000", 
160 => x"71fc0608", 
161 => x"0b0b0bb4", 
162 => x"94738306", 
163 => x"10100508", 
164 => x"060b0b0b", 
165 => x"88a20400", 
166 => x"00000000", 
167 => x"00000000", 
168 => x"88088c08", 
169 => x"90087575", 
170 => x"0b0b0bb1", 
171 => x"bd2d5050", 
172 => x"88085690", 
173 => x"0c8c0c88", 
174 => x"0c510400", 
175 => x"00000000", 
176 => x"88088c08", 
177 => x"90087575", 
178 => x"0b0b0bb1", 
179 => x"f82d5050", 
180 => x"88085690", 
181 => x"0c8c0c88", 
182 => x"0c510400", 
183 => x"00000000", 
184 => x"72097081", 
185 => x"0509060a", 
186 => x"8106ff05", 
187 => x"70547106", 
188 => x"73097274", 
189 => x"05ff0506", 
190 => x"07515151", 
191 => x"04000000", 
192 => x"72097081", 
193 => x"0509060a", 
194 => x"098106ff", 
195 => x"05705471", 
196 => x"06730972", 
197 => x"7405ff05", 
198 => x"06075151", 
199 => x"51040000", 
200 => x"05ff0504", 
201 => x"00000000", 
202 => x"00000000", 
203 => x"00000000", 
204 => x"00000000", 
205 => x"00000000", 
206 => x"00000000", 
207 => x"00000000", 
208 => x"04000000", 
209 => x"00000000", 
210 => x"00000000", 
211 => x"00000000", 
212 => x"00000000", 
213 => x"00000000", 
214 => x"00000000", 
215 => x"00000000", 
216 => x"71810552", 
217 => x"04000000", 
218 => x"00000000", 
219 => x"00000000", 
220 => x"00000000", 
221 => x"00000000", 
222 => x"00000000", 
223 => x"00000000", 
224 => x"04000000", 
225 => x"00000000", 
226 => x"00000000", 
227 => x"00000000", 
228 => x"00000000", 
229 => x"00000000", 
230 => x"00000000", 
231 => x"00000000", 
232 => x"02840572", 
233 => x"10100552", 
234 => x"04000000", 
235 => x"00000000", 
236 => x"00000000", 
237 => x"00000000", 
238 => x"00000000", 
239 => x"00000000", 
240 => x"00000000", 
241 => x"00000000", 
242 => x"00000000", 
243 => x"00000000", 
244 => x"00000000", 
245 => x"00000000", 
246 => x"00000000", 
247 => x"00000000", 
248 => x"717105ff", 
249 => x"05715351", 
250 => x"020d0400", 
251 => x"00000000", 
252 => x"00000000", 
253 => x"00000000", 
254 => x"00000000", 
255 => x"00000000", 
256 => x"10101010", 
257 => x"10101010", 
258 => x"10101010", 
259 => x"10101010", 
260 => x"10101010", 
261 => x"10101010", 
262 => x"10101010", 
263 => x"10101053", 
264 => x"51047381", 
265 => x"ff067383", 
266 => x"06098105", 
267 => x"83051010", 
268 => x"102b0772", 
269 => x"fc060c51", 
270 => x"51047272", 
271 => x"80728106", 
272 => x"ff050972", 
273 => x"06057110", 
274 => x"52720a10", 
275 => x"0a5372ed", 
276 => x"38515153", 
277 => x"51040000", 
278 => x"80040088", 
279 => x"da040400", 
280 => x"00000004", 
281 => x"5eb8c870", 
282 => x"80c1c427", 
283 => x"8b388071", 
284 => x"70840553", 
285 => x"0c88e704", 
286 => x"88da5196", 
287 => x"d90402f8", 
288 => x"050d7352", 
289 => x"c0087088", 
290 => x"2a708106", 
291 => x"51515170", 
292 => x"802ef138", 
293 => x"71c00c71", 
294 => x"880c0288", 
295 => x"050d0402", 
296 => x"f0050d75", 
297 => x"537284e0", 
298 => x"2d7081ff", 
299 => x"06525270", 
300 => x"802ea238", 
301 => x"7181ff06", 
302 => x"81145452", 
303 => x"c0087088", 
304 => x"2a708106", 
305 => x"51515170", 
306 => x"802ef138", 
307 => x"71c00c81", 
308 => x"145489a5", 
309 => x"0473880c", 
310 => x"0290050d", 
311 => x"0402f805", 
312 => x"0dc00870", 
313 => x"892a7081", 
314 => x"06515252", 
315 => x"70802ef1", 
316 => x"387181ff", 
317 => x"06880c02", 
318 => x"88050d04", 
319 => x"02f4050d", 
320 => x"94f32d88", 
321 => x"08b8b408", 
322 => x"055394f3", 
323 => x"2d728808", 
324 => x"27863880", 
325 => x"518ab104", 
326 => x"c0087089", 
327 => x"2a708106", 
328 => x"51525270", 
329 => x"802ee338", 
330 => x"74517171", 
331 => x"85802d81", 
332 => x"5170880c", 
333 => x"028c050d", 
334 => x"0402f405", 
335 => x"0dd45281", 
336 => x"ff720c71", 
337 => x"085381ff", 
338 => x"720c7288", 
339 => x"2b83fe80", 
340 => x"06720870", 
341 => x"81ff0651", 
342 => x"525381ff", 
343 => x"720c7271", 
344 => x"07882b72", 
345 => x"087081ff", 
346 => x"06515253", 
347 => x"81ff720c", 
348 => x"72710788", 
349 => x"2b720870", 
350 => x"81ff0672", 
351 => x"07880c52", 
352 => x"53028c05", 
353 => x"0d0402f4", 
354 => x"050d7476", 
355 => x"7181ff06", 
356 => x"d40c5353", 
357 => x"bcec0885", 
358 => x"3871892b", 
359 => x"5271982a", 
360 => x"d40c7190", 
361 => x"2a7081ff", 
362 => x"06d40c51", 
363 => x"71882a70", 
364 => x"81ff06d4", 
365 => x"0c517181", 
366 => x"ff06d40c", 
367 => x"72902a70", 
368 => x"81ff06d4", 
369 => x"0c51d408", 
370 => x"7081ff06", 
371 => x"515182b8", 
372 => x"bf527081", 
373 => x"ff2e0981", 
374 => x"06943881", 
375 => x"ff0bd40c", 
376 => x"d4087081", 
377 => x"ff06ff14", 
378 => x"54515171", 
379 => x"e5387088", 
380 => x"0c028c05", 
381 => x"0d0402fc", 
382 => x"050d81c7", 
383 => x"5181ff0b", 
384 => x"d40cff11", 
385 => x"51708025", 
386 => x"f4380284", 
387 => x"050d0402", 
388 => x"f0050d8b", 
389 => x"f62d819c", 
390 => x"9f538052", 
391 => x"87fc80f7", 
392 => x"518b862d", 
393 => x"88085488", 
394 => x"08812e09", 
395 => x"8106a238", 
396 => x"81ff0bd4", 
397 => x"0c820a52", 
398 => x"849c80e9", 
399 => x"518b862d", 
400 => x"88088b38", 
401 => x"81ff0bd4", 
402 => x"0c73538c", 
403 => x"d7048bf6", 
404 => x"2dff1353", 
405 => x"72c43872", 
406 => x"880c0290", 
407 => x"050d0402", 
408 => x"f4050d81", 
409 => x"ff0bd40c", 
410 => x"93538052", 
411 => x"87fc80c1", 
412 => x"518b862d", 
413 => x"88088b38", 
414 => x"81ff0bd4", 
415 => x"0c81538d", 
416 => x"8b048bf6", 
417 => x"2dff1353", 
418 => x"72e03872", 
419 => x"880c028c", 
420 => x"050d0402", 
421 => x"f0050d8b", 
422 => x"f62d83aa", 
423 => x"52849c80", 
424 => x"c8518b86", 
425 => x"2d880881", 
426 => x"2e098106", 
427 => x"91388ab9", 
428 => x"2d880883", 
429 => x"ffff0653", 
430 => x"7283aa2e", 
431 => x"91388cdf", 
432 => x"2d8dc904", 
433 => x"81548eaa", 
434 => x"0480548e", 
435 => x"aa0481ff", 
436 => x"0bd40cb1", 
437 => x"538c8f2d", 
438 => x"8808802e", 
439 => x"be388052", 
440 => x"87fc80fa", 
441 => x"518b862d", 
442 => x"8808b038", 
443 => x"81ff0bd4", 
444 => x"0cd40853", 
445 => x"81ff0bd4", 
446 => x"0c81ff0b", 
447 => x"d40c81ff", 
448 => x"0bd40c81", 
449 => x"ff0bd40c", 
450 => x"72862a70", 
451 => x"81068808", 
452 => x"56515372", 
453 => x"802e9338", 
454 => x"8dc40472", 
455 => x"822effa9", 
456 => x"38ff1353", 
457 => x"72ffae38", 
458 => x"72547388", 
459 => x"0c029005", 
460 => x"0d0402e8", 
461 => x"050d7856", 
462 => x"81ff0bd4", 
463 => x"0cd00870", 
464 => x"8f2a7081", 
465 => x"06515153", 
466 => x"72f33882", 
467 => x"810bd00c", 
468 => x"81ff0bd4", 
469 => x"0c775287", 
470 => x"fc80d851", 
471 => x"8b862d81", 
472 => x"53880880", 
473 => x"f93881ff", 
474 => x"0bd40c81", 
475 => x"fe0bd40c", 
476 => x"80ff5575", 
477 => x"70840557", 
478 => x"0870982a", 
479 => x"d40c7090", 
480 => x"2c7081ff", 
481 => x"06d40c54", 
482 => x"70882c70", 
483 => x"81ff06d4", 
484 => x"0c547081", 
485 => x"ff06d40c", 
486 => x"54ff1555", 
487 => x"748025d3", 
488 => x"3881ff0b", 
489 => x"d40c81ff", 
490 => x"0bd40c81", 
491 => x"ff0bd40c", 
492 => x"868da054", 
493 => x"81ff0bd4", 
494 => x"0cd40881", 
495 => x"ff065574", 
496 => x"8738ff14", 
497 => x"5473ed38", 
498 => x"81ff0bd4", 
499 => x"0cd00870", 
500 => x"8f2a7081", 
501 => x"06515153", 
502 => x"72f33872", 
503 => x"d00c7288", 
504 => x"0c029805", 
505 => x"0d0402ec", 
506 => x"050d7678", 
507 => x"53548055", 
508 => x"80dbc6df", 
509 => x"5381ff0b", 
510 => x"d40cd408", 
511 => x"7081ff06", 
512 => x"51517081", 
513 => x"fe2e0981", 
514 => x"0680cc38", 
515 => x"800bbd90", 
516 => x"0c837225", 
517 => x"9b388ab9", 
518 => x"2d880874", 
519 => x"70840556", 
520 => x"0cbd9008", 
521 => x"880805bd", 
522 => x"900cfc12", 
523 => x"52909104", 
524 => x"8072259e", 
525 => x"3881ff0b", 
526 => x"d40cff74", 
527 => x"70810556", 
528 => x"85802dbd", 
529 => x"900881ff", 
530 => x"05bd900c", 
531 => x"ff125290", 
532 => x"b0048155", 
533 => x"90de04ff", 
534 => x"135372ff", 
535 => x"983881ff", 
536 => x"0bd40c74", 
537 => x"880c0294", 
538 => x"050d0402", 
539 => x"e8050d80", 
540 => x"5287fc80", 
541 => x"c9518b86", 
542 => x"2d9252bc", 
543 => x"fc518fe6", 
544 => x"2dbcfc0b", 
545 => x"84e02d81", 
546 => x"c0065372", 
547 => x"80c02e09", 
548 => x"8106b038", 
549 => x"bd830b84", 
550 => x"e02dbd84", 
551 => x"0b84e02d", 
552 => x"71902b71", 
553 => x"882b07bd", 
554 => x"850b84e0", 
555 => x"2d7181ff", 
556 => x"fe800607", 
557 => x"70888029", 
558 => x"88800551", 
559 => x"51555755", 
560 => x"92ad04bd", 
561 => x"850b84e0", 
562 => x"2d701086", 
563 => x"06bd860b", 
564 => x"84e02d70", 
565 => x"872a7207", 
566 => x"bd810b84", 
567 => x"e02d8f06", 
568 => x"bd820b84", 
569 => x"e02d708a", 
570 => x"2b988006", 
571 => x"bd830b84", 
572 => x"e02d7082", 
573 => x"2b7207bd", 
574 => x"840b84e0", 
575 => x"2d70862a", 
576 => x"72078218", 
577 => x"81782b81", 
578 => x"1381732b", 
579 => x"71295153", 
580 => x"58585252", 
581 => x"52525953", 
582 => x"54525855", 
583 => x"55848075", 
584 => x"258b3872", 
585 => x"1075812c", 
586 => x"5653929d", 
587 => x"0472880c", 
588 => x"0298050d", 
589 => x"0402f005", 
590 => x"0d810bbc", 
591 => x"ec0c8754", 
592 => x"d008708f", 
593 => x"2a708106", 
594 => x"51515372", 
595 => x"f33872d0", 
596 => x"0c8bf62d", 
597 => x"d008708f", 
598 => x"2a708106", 
599 => x"51515372", 
600 => x"f338810b", 
601 => x"d00c7252", 
602 => x"84d480c0", 
603 => x"518b862d", 
604 => x"8808812e", 
605 => x"8e387382", 
606 => x"2e80c338", 
607 => x"ff145473", 
608 => x"ffbe388d", 
609 => x"932d8808", 
610 => x"bcec0c88", 
611 => x"088b3881", 
612 => x"5287fc80", 
613 => x"d0518b86", 
614 => x"2d81ff0b", 
615 => x"d40c90eb", 
616 => x"2d8808bc", 
617 => x"f00cd008", 
618 => x"708f2a70", 
619 => x"81065151", 
620 => x"5372f338", 
621 => x"72d00c81", 
622 => x"ff0bd40c", 
623 => x"81537288", 
624 => x"0c029005", 
625 => x"0d0402f0", 
626 => x"050d8054", 
627 => x"81ff0bd4", 
628 => x"0cd00870", 
629 => x"8f2a7081", 
630 => x"06515153", 
631 => x"72f33882", 
632 => x"810bd00c", 
633 => x"81ff0bd4", 
634 => x"0c755287", 
635 => x"fc80d151", 
636 => x"8b862d88", 
637 => x"089d3884", 
638 => x"80527651", 
639 => x"8fe62d88", 
640 => x"0854d008", 
641 => x"708f2a70", 
642 => x"81065151", 
643 => x"5372f338", 
644 => x"72d00c73", 
645 => x"880c0290", 
646 => x"050d0402", 
647 => x"f4050d74", 
648 => x"70882a83", 
649 => x"fe800670", 
650 => x"72982a07", 
651 => x"72882b87", 
652 => x"fc808006", 
653 => x"71077398", 
654 => x"2b07880c", 
655 => x"51535102", 
656 => x"8c050d04", 
657 => x"02f8050d", 
658 => x"028e0584", 
659 => x"e02d7488", 
660 => x"2b077083", 
661 => x"ffff0688", 
662 => x"0c510288", 
663 => x"050d0402", 
664 => x"f8050d73", 
665 => x"70902b71", 
666 => x"902a0788", 
667 => x"0c520288", 
668 => x"050d04c8", 
669 => x"08880c04", 
670 => x"810b880c", 
671 => x"0402dc05", 
672 => x"0d7a5202", 
673 => x"a405ec05", 
674 => x"51a5b92d", 
675 => x"8808802e", 
676 => x"80f73876", 
677 => x"0b0b0bbc", 
678 => x"d80c0b0b", 
679 => x"0bb8c852", 
680 => x"02900570", 
681 => x"5254a7bb", 
682 => x"2d800b0b", 
683 => x"0b0bbcd4", 
684 => x"0c0b0b0b", 
685 => x"bcd80880", 
686 => x"2ebf380b", 
687 => x"0b0bbcd4", 
688 => x"080b0b0b", 
689 => x"b8c80570", 
690 => x"84e02d52", 
691 => x"5388fe2d", 
692 => x"0b0b0bbc", 
693 => x"d808ff05", 
694 => x"0b0b0bbc", 
695 => x"d80c0b0b", 
696 => x"0bbcd408", 
697 => x"81050b0b", 
698 => x"0bbcd40c", 
699 => x"83ff0b0b", 
700 => x"0b0bbcd4", 
701 => x"0825ffb9", 
702 => x"38815273", 
703 => x"51a6f02d", 
704 => x"0b0b0bbc", 
705 => x"d808ff92", 
706 => x"3802a405", 
707 => x"0d0402fc", 
708 => x"050d94f3", 
709 => x"2d880813", 
710 => x"5194f32d", 
711 => x"70880827", 
712 => x"f8380284", 
713 => x"050d0402", 
714 => x"f4050d74", 
715 => x"53807325", 
716 => x"9f387252", 
717 => x"810bffa0", 
718 => x"0c81fa51", 
719 => x"968e2d80", 
720 => x"0bffa00c", 
721 => x"81fa5196", 
722 => x"8e2dff12", 
723 => x"5271e538", 
724 => x"87e85196", 
725 => x"8e2d96ad", 
726 => x"0402dc05", 
727 => x"0d817059", 
728 => x"5792b52d", 
729 => x"9ce52db4", 
730 => x"a451ad93", 
731 => x"2d83f40b", 
732 => x"b8b40c02", 
733 => x"a405fc05", 
734 => x"5189fc2d", 
735 => x"88089f38", 
736 => x"ffa80870", 
737 => x"78068106", 
738 => x"51547380", 
739 => x"2ee53888", 
740 => x"085787e8", 
741 => x"51968e2d", 
742 => x"b788519b", 
743 => x"ac0402a0", 
744 => x"0584e02d", 
745 => x"51b3f12d", 
746 => x"8808ffbf", 
747 => x"05547393", 
748 => x"26c13873", 
749 => x"8429b4b4", 
750 => x"05547308", 
751 => x"0489dd2d", 
752 => x"88080b0b", 
753 => x"0bbcc80b", 
754 => x"85802d80", 
755 => x"0b880881", 
756 => x"ff065555", 
757 => x"73752e83", 
758 => x"38815574", 
759 => x"ffa40c96", 
760 => x"f304800b", 
761 => x"0b0b0bbc", 
762 => x"d40c0b0b", 
763 => x"0bbcd408", 
764 => x"0b0b0bbc", 
765 => x"c8055489", 
766 => x"dd2d8808", 
767 => x"7485802d", 
768 => x"0b0b0bbc", 
769 => x"d4088105", 
770 => x"0b0b0bbc", 
771 => x"d40c8a0b", 
772 => x"0b0b0bbc", 
773 => x"d40825d2", 
774 => x"38800b0b", 
775 => x"0b0bbcd3", 
776 => x"0b85802d", 
777 => x"8b53b794", 
778 => x"520b0b0b", 
779 => x"bcc8519c", 
780 => x"a32d8808", 
781 => x"95387780", 
782 => x"2e873888", 
783 => x"085896f3", 
784 => x"04880851", 
785 => x"aeaa2d96", 
786 => x"f3040b0b", 
787 => x"0bbcc851", 
788 => x"ad932d96", 
789 => x"f30494f8", 
790 => x"528151a3", 
791 => x"8f2d8808", 
792 => x"bd940cbd", 
793 => x"94088b11", 
794 => x"84e02d70", 
795 => x"842a7081", 
796 => x"06515657", 
797 => x"5573802e", 
798 => x"80cc388b", 
799 => x"53b7a052", 
800 => x"74519ca3", 
801 => x"2d880880", 
802 => x"2e81a438", 
803 => x"800b0b0b", 
804 => x"0bbcd40c", 
805 => x"0b0b0bbc", 
806 => x"d408bd94", 
807 => x"08057084", 
808 => x"e02d5254", 
809 => x"88fe2d0b", 
810 => x"0b0bbcd4", 
811 => x"0881050b", 
812 => x"0b0bbcd4", 
813 => x"0c8a0b0b", 
814 => x"0b0bbcd4", 
815 => x"0825d538", 
816 => x"80d1519a", 
817 => x"a7047598", 
818 => x"06547380", 
819 => x"e2388353", 
820 => x"b7905288", 
821 => x"15519ca3", 
822 => x"2d880880", 
823 => x"2e933883", 
824 => x"53b7ac52", 
825 => x"bd940888", 
826 => x"05519ca3", 
827 => x"2d8808bf", 
828 => x"38730b0b", 
829 => x"0bbcd40c", 
830 => x"0b0b0bbc", 
831 => x"d408bd94", 
832 => x"08057084", 
833 => x"e02d5254", 
834 => x"88fe2d0b", 
835 => x"0b0bbcd4", 
836 => x"0881050b", 
837 => x"0b0bbcd4", 
838 => x"0c8a0b0b", 
839 => x"0b0bbcd4", 
840 => x"0825d538", 
841 => x"80f15188", 
842 => x"fe2d8051", 
843 => x"88fe2d94", 
844 => x"f8528051", 
845 => x"a38f2d88", 
846 => x"08bd940c", 
847 => x"8808fea3", 
848 => x"3881ff51", 
849 => x"9c9d0489", 
850 => x"dd2d8808", 
851 => x"0b0b0bbc", 
852 => x"c80b8580", 
853 => x"2d880881", 
854 => x"ff06519c", 
855 => x"9d04800b", 
856 => x"0b0b0bbc", 
857 => x"d40c0b0b", 
858 => x"0bbcd408", 
859 => x"0b0b0bbc", 
860 => x"c8055489", 
861 => x"dd2d8808", 
862 => x"7485802d", 
863 => x"0b0b0bbc", 
864 => x"d4088105", 
865 => x"0b0b0bbc", 
866 => x"d40c8a0b", 
867 => x"0b0b0bbc", 
868 => x"d40825d2", 
869 => x"38800b0b", 
870 => x"0b0bbcd3", 
871 => x"0b85802d", 
872 => x"87e85196", 
873 => x"8e2d0b0b", 
874 => x"0bbcc851", 
875 => x"94fd2d96", 
876 => x"f30489dd", 
877 => x"2d88080b", 
878 => x"0b0bbcc8", 
879 => x"0b85802d", 
880 => x"800b8808", 
881 => x"81ff0655", 
882 => x"5573752e", 
883 => x"83388155", 
884 => x"74ffa00c", 
885 => x"96f30492", 
886 => x"519c9d04", 
887 => x"815796f3", 
888 => x"04b7b051", 
889 => x"899f2d80", 
890 => x"519c9d04", 
891 => x"805796f3", 
892 => x"04ab519c", 
893 => x"9d0482ac", 
894 => x"51968e2d", 
895 => x"825188fe", 
896 => x"2d80c751", 
897 => x"88fe2d91", 
898 => x"5188fe2d", 
899 => x"825188fe", 
900 => x"2d835188", 
901 => x"fe2d8851", 
902 => x"88fe2d89", 
903 => x"5188fe2d", 
904 => x"96f30402", 
905 => x"e8050d77", 
906 => x"797b5855", 
907 => x"55805372", 
908 => x"7625a338", 
909 => x"74708105", 
910 => x"5684e02d", 
911 => x"74708105", 
912 => x"5684e02d", 
913 => x"52527171", 
914 => x"2e863881", 
915 => x"519cd804", 
916 => x"8113539c", 
917 => x"af048051", 
918 => x"70880c02", 
919 => x"98050d04", 
920 => x"810b880c", 
921 => x"0402d805", 
922 => x"0d800b80", 
923 => x"c1b00cbd", 
924 => x"a0528051", 
925 => x"93c62d88", 
926 => x"08558808", 
927 => x"802e858e", 
928 => x"38805688", 
929 => x"53b8b808", 
930 => x"52bdd651", 
931 => x"b3a52d88", 
932 => x"08810509", 
933 => x"70880807", 
934 => x"9f2a5154", 
935 => x"8853b8bc", 
936 => x"0852bdf2", 
937 => x"51b3a52d", 
938 => x"8808762e", 
939 => x"80ff3873", 
940 => x"762e80f9", 
941 => x"3880c0e6", 
942 => x"0b84e02d", 
943 => x"80c0e70b", 
944 => x"84e02d71", 
945 => x"982b7190", 
946 => x"2b0780c0", 
947 => x"e80b84e0", 
948 => x"2d70882b", 
949 => x"720780c0", 
950 => x"e90b84e0", 
951 => x"2d710780", 
952 => x"c19e0b84", 
953 => x"e02d80c1", 
954 => x"9f0b84e0", 
955 => x"2d71882b", 
956 => x"07535f54", 
957 => x"525a5657", 
958 => x"557381ab", 
959 => x"aa2e0981", 
960 => x"068c3875", 
961 => x"51949b2d", 
962 => x"8808569e", 
963 => x"9b048055", 
964 => x"7382d4d5", 
965 => x"2e098106", 
966 => x"83f438bd", 
967 => x"a0527551", 
968 => x"93c62d88", 
969 => x"08558808", 
970 => x"802e83e2", 
971 => x"388853b8", 
972 => x"bc0852bd", 
973 => x"f251b3a5", 
974 => x"2d88088a", 
975 => x"38810b80", 
976 => x"c1b00c9e", 
977 => x"de048853", 
978 => x"b8b80852", 
979 => x"bdd651b3", 
980 => x"a52d8055", 
981 => x"8808752e", 
982 => x"09810683", 
983 => x"b13880c1", 
984 => x"9e0b84e0", 
985 => x"2d547380", 
986 => x"d52e0981", 
987 => x"0680cb38", 
988 => x"80c19f0b", 
989 => x"84e02d54", 
990 => x"7381aa2e", 
991 => x"098106ba", 
992 => x"38800bbd", 
993 => x"a00b84e0", 
994 => x"2d565474", 
995 => x"81e92e83", 
996 => x"38815474", 
997 => x"81eb2e8c", 
998 => x"38805573", 
999 => x"752e0981", 
1000 => x"0682eb38", 
1001 => x"bdab0b84", 
1002 => x"e02d5574", 
1003 => x"8d38bdac", 
1004 => x"0b84e02d", 
1005 => x"5473822e", 
1006 => x"86388055", 
1007 => x"a28e04bd", 
1008 => x"ad0b84e0", 
1009 => x"2d7080c1", 
1010 => x"bc0cff11", 
1011 => x"80c1ac0c", 
1012 => x"bdae0b84", 
1013 => x"e02dbdaf", 
1014 => x"0b84e02d", 
1015 => x"5a770579", 
1016 => x"82802905", 
1017 => x"7080c1a4", 
1018 => x"0cbdb00b", 
1019 => x"84e02d80", 
1020 => x"c1b0085b", 
1021 => x"5b575777", 
1022 => x"802e8199", 
1023 => x"388853b8", 
1024 => x"bc0852bd", 
1025 => x"f251b3a5", 
1026 => x"2d880882", 
1027 => x"81387684", 
1028 => x"2b80c1a0", 
1029 => x"0c7680c1", 
1030 => x"b80cbdc5", 
1031 => x"0b84e02d", 
1032 => x"bdc40b84", 
1033 => x"e02d7182", 
1034 => x"802905bd", 
1035 => x"c60b84e0", 
1036 => x"2d708480", 
1037 => x"802912bd", 
1038 => x"c70b84e0", 
1039 => x"2d527181", 
1040 => x"800a2905", 
1041 => x"7c71291a", 
1042 => x"7080c1c0", 
1043 => x"0cbdcd0b", 
1044 => x"84e02dbd", 
1045 => x"cc0b84e0", 
1046 => x"2d718280", 
1047 => x"2905bdce", 
1048 => x"0b84e02d", 
1049 => x"70848080", 
1050 => x"2912bdcf", 
1051 => x"0b84e02d", 
1052 => x"70982b81", 
1053 => x"f00a0672", 
1054 => x"0570bd9c", 
1055 => x"0cfe1162", 
1056 => x"29770580", 
1057 => x"c1a80c52", 
1058 => x"42525555", 
1059 => x"525a5852", 
1060 => x"555aa1e3", 
1061 => x"04bdb20b", 
1062 => x"84e02dbd", 
1063 => x"b10b84e0", 
1064 => x"2d718280", 
1065 => x"29057080", 
1066 => x"c1a00c70", 
1067 => x"a02983ff", 
1068 => x"0570892a", 
1069 => x"7080c1b8", 
1070 => x"0cbdb70b", 
1071 => x"84e02dbd", 
1072 => x"b60b84e0", 
1073 => x"2d718280", 
1074 => x"29057e71", 
1075 => x"291c7080", 
1076 => x"c1a80c7e", 
1077 => x"bd9c0c73", 
1078 => x"0580c1c0", 
1079 => x"0c5a5b51", 
1080 => x"51555abd", 
1081 => x"9c08bd98", 
1082 => x"0c80c1a8", 
1083 => x"0880c1b4", 
1084 => x"0c77802e", 
1085 => x"8b3880c1", 
1086 => x"bc08842b", 
1087 => x"54a28704", 
1088 => x"80c1b808", 
1089 => x"842b5473", 
1090 => x"80c1a00c", 
1091 => x"81557488", 
1092 => x"0c02a805", 
1093 => x"0d0402ec", 
1094 => x"050d7670", 
1095 => x"872a7180", 
1096 => x"ff065754", 
1097 => x"5480c1b0", 
1098 => x"088a3873", 
1099 => x"882a7481", 
1100 => x"ff065653", 
1101 => x"80c1a408", 
1102 => x"1353b8c0", 
1103 => x"08732e96", 
1104 => x"3872b8c0", 
1105 => x"0cbda052", 
1106 => x"725193c6", 
1107 => x"2d880853", 
1108 => x"8808802e", 
1109 => x"b23880c1", 
1110 => x"b008802e", 
1111 => x"97387484", 
1112 => x"29bda005", 
1113 => x"70085253", 
1114 => x"949b2d88", 
1115 => x"08f00a06", 
1116 => x"55a38504", 
1117 => x"7410bda0", 
1118 => x"057080c0", 
1119 => x"2d525394", 
1120 => x"c42d8808", 
1121 => x"55745372", 
1122 => x"880c0294", 
1123 => x"050d0402", 
1124 => x"e0050d7a", 
1125 => x"5879802e", 
1126 => x"9338800b", 
1127 => x"bce80c80", 
1128 => x"c1b408bc", 
1129 => x"e00cbd98", 
1130 => x"08bce40c", 
1131 => x"bce80853", 
1132 => x"7280c1a0", 
1133 => x"08278197", 
1134 => x"38728f06", 
1135 => x"5372a238", 
1136 => x"bce008b8", 
1137 => x"c00cbda0", 
1138 => x"52bce008", 
1139 => x"51bce008", 
1140 => x"8105bce0", 
1141 => x"0c93c62d", 
1142 => x"bda00bbc", 
1143 => x"dc0ca3e9", 
1144 => x"04bcdc08", 
1145 => x"a005bcdc", 
1146 => x"0cbce808", 
1147 => x"8105bce8", 
1148 => x"0c800bbc", 
1149 => x"dc087084", 
1150 => x"e02d5557", 
1151 => x"5472742e", 
1152 => x"83388154", 
1153 => x"7281e52e", 
1154 => x"ffa23881", 
1155 => x"70750654", 
1156 => x"5772802e", 
1157 => x"ff96388b", 
1158 => x"1684e02d", 
1159 => x"70832a78", 
1160 => x"06565474", 
1161 => x"ff863873", 
1162 => x"842a7078", 
1163 => x"06765651", 
1164 => x"53778338", 
1165 => x"76547274", 
1166 => x"0753728c", 
1167 => x"38755177", 
1168 => x"2d880880", 
1169 => x"2efee538", 
1170 => x"bcdc0853", 
1171 => x"a5b10480", 
1172 => x"c1b4088a", 
1173 => x"3880c1b0", 
1174 => x"08802e80", 
1175 => x"d238bce4", 
1176 => x"0851a296", 
1177 => x"2d8808bc", 
1178 => x"e40c80c1", 
1179 => x"b008802e", 
1180 => x"96388808", 
1181 => x"80ffffff", 
1182 => x"f8065372", 
1183 => x"80ffffff", 
1184 => x"f82eac38", 
1185 => x"a5950488", 
1186 => x"0883fff8", 
1187 => x"06537283", 
1188 => x"fff82e9b", 
1189 => x"38bce408", 
1190 => x"fe0580c1", 
1191 => x"bc082980", 
1192 => x"c1c00805", 
1193 => x"bce00c80", 
1194 => x"0bbce80c", 
1195 => x"a3ac0480", 
1196 => x"5372880c", 
1197 => x"02a0050d", 
1198 => x"0402e405", 
1199 => x"0d787a56", 
1200 => x"57807055", 
1201 => x"5676762e", 
1202 => x"819e3875", 
1203 => x"88180c74", 
1204 => x"762e8192", 
1205 => x"387484e0", 
1206 => x"2d547376", 
1207 => x"2e818738", 
1208 => x"9ce05281", 
1209 => x"51a38f2d", 
1210 => x"a5fb048b", 
1211 => x"53745288", 
1212 => x"08519ca3", 
1213 => x"2d880880", 
1214 => x"2e93389c", 
1215 => x"e0528051", 
1216 => x"a38f2d88", 
1217 => x"08568808", 
1218 => x"e238a6e6", 
1219 => x"0475802e", 
1220 => x"80d4389c", 
1221 => x"16085194", 
1222 => x"9b2d8808", 
1223 => x"88180c9a", 
1224 => x"1680c02d", 
1225 => x"5194c42d", 
1226 => x"88088808", 
1227 => x"84190c88", 
1228 => x"08555580", 
1229 => x"c1b00880", 
1230 => x"2e973894", 
1231 => x"1680c02d", 
1232 => x"5194c42d", 
1233 => x"8808902b", 
1234 => x"83fff00a", 
1235 => x"06701651", 
1236 => x"54738418", 
1237 => x"0c80770c", 
1238 => x"738c180c", 
1239 => x"800b9018", 
1240 => x"0c8154a6", 
1241 => x"e8047554", 
1242 => x"73880c02", 
1243 => x"9c050d04", 
1244 => x"02ec050d", 
1245 => x"76785654", 
1246 => x"73802eba", 
1247 => x"38881408", 
1248 => x"802eb338", 
1249 => x"73087016", 
1250 => x"565280c1", 
1251 => x"ac080972", 
1252 => x"76320652", 
1253 => x"71802e9b", 
1254 => x"38841408", 
1255 => x"51a2962d", 
1256 => x"88088415", 
1257 => x"0c730880", 
1258 => x"c1bc0805", 
1259 => x"70750c52", 
1260 => x"a78a0474", 
1261 => x"740c0294", 
1262 => x"050d0402", 
1263 => x"f0050d75", 
1264 => x"5473802e", 
1265 => x"86388814", 
1266 => x"08863880", 
1267 => x"53a7fd04", 
1268 => x"841408fe", 
1269 => x"0580c1bc", 
1270 => x"082980c1", 
1271 => x"c0081175", 
1272 => x"0880c1ac", 
1273 => x"08060570", 
1274 => x"b8c00c78", 
1275 => x"54525393", 
1276 => x"c62d8808", 
1277 => x"53880880", 
1278 => x"2e833881", 
1279 => x"5372880c", 
1280 => x"0290050d", 
1281 => x"0402f005", 
1282 => x"0d755473", 
1283 => x"802e8638", 
1284 => x"88140886", 
1285 => x"388053a8", 
1286 => x"c7048414", 
1287 => x"08fe0580", 
1288 => x"c1bc0829", 
1289 => x"80c1c008", 
1290 => x"11750880", 
1291 => x"c1ac0806", 
1292 => x"0570b8c0", 
1293 => x"0c785452", 
1294 => x"538eb22d", 
1295 => x"88085388", 
1296 => x"08802e83", 
1297 => x"38815372", 
1298 => x"880c0290", 
1299 => x"050d0402", 
1300 => x"e4050d78", 
1301 => x"7a705957", 
1302 => x"5473802e", 
1303 => x"80cb3888", 
1304 => x"1408802e", 
1305 => x"80c33880", 
1306 => x"c1ac0809", 
1307 => x"90150870", 
1308 => x"72065256", 
1309 => x"53757327", 
1310 => x"92388074", 
1311 => x"0c800b90", 
1312 => x"150c8c14", 
1313 => x"0884150c", 
1314 => x"a9940474", 
1315 => x"fc800676", 
1316 => x"71315853", 
1317 => x"76892a52", 
1318 => x"7351a6f0", 
1319 => x"2dbda052", 
1320 => x"7351a7bb", 
1321 => x"2d759015", 
1322 => x"0c029c05", 
1323 => x"0d0402e0", 
1324 => x"050d797b", 
1325 => x"7d575858", 
1326 => x"77802e88", 
1327 => x"38881808", 
1328 => x"54738638", 
1329 => x"8053aafe", 
1330 => x"04901808", 
1331 => x"70165456", 
1332 => x"73732785", 
1333 => x"38737631", 
1334 => x"55805372", 
1335 => x"7525819e", 
1336 => x"387583ff", 
1337 => x"06547373", 
1338 => x"2ebc3884", 
1339 => x"807431bd", 
1340 => x"a0155553", 
1341 => x"74732583", 
1342 => x"38745372", 
1343 => x"1690190c", 
1344 => x"74733155", 
1345 => x"ff135372", 
1346 => x"ff2e9438", 
1347 => x"73708105", 
1348 => x"5584e02d", 
1349 => x"77708105", 
1350 => x"5985802d", 
1351 => x"aa840481", 
1352 => x"527751a6", 
1353 => x"f02d8153", 
1354 => x"80752580", 
1355 => x"d13883ff", 
1356 => x"75259c38", 
1357 => x"76527751", 
1358 => x"a7bb2d84", 
1359 => x"80179019", 
1360 => x"08848005", 
1361 => x"901a0cfc", 
1362 => x"80165657", 
1363 => x"aa9f04bd", 
1364 => x"a0527751", 
1365 => x"a7bb2dbd", 
1366 => x"a00b9019", 
1367 => x"0816901a", 
1368 => x"0c54ff15", 
1369 => x"5574ff2e", 
1370 => x"ffb53873", 
1371 => x"70810555", 
1372 => x"84e02d77", 
1373 => x"70810559", 
1374 => x"85802daa", 
1375 => x"e2047288", 
1376 => x"0c02a005", 
1377 => x"0d0402ec", 
1378 => x"050d7654", 
1379 => x"73802e86", 
1380 => x"38881408", 
1381 => x"8638ff53", 
1382 => x"abda0490", 
1383 => x"14087083", 
1384 => x"ff065455", 
1385 => x"72953874", 
1386 => x"802e8838", 
1387 => x"81527351", 
1388 => x"a6f02dbd", 
1389 => x"a0527351", 
1390 => x"a7bb2d90", 
1391 => x"140855ff", 
1392 => x"53748815", 
1393 => x"08279338", 
1394 => x"7483ff06", 
1395 => x"bda00570", 
1396 => x"84e02d81", 
1397 => x"1790170c", 
1398 => x"51537288", 
1399 => x"0c029405", 
1400 => x"0d0402d8", 
1401 => x"050d7c7c", 
1402 => x"53029805", 
1403 => x"70535653", 
1404 => x"a5b92d88", 
1405 => x"08548808", 
1406 => x"802eb438", 
1407 => x"80547774", 
1408 => x"2eab3872", 
1409 => x"527451a7", 
1410 => x"bb2d8808", 
1411 => x"802e9838", 
1412 => x"81527451", 
1413 => x"a6f02d84", 
1414 => x"80138480", 
1415 => x"15555377", 
1416 => x"7426e038", 
1417 => x"acad0488", 
1418 => x"0854acaf", 
1419 => x"04815473", 
1420 => x"880c02a8", 
1421 => x"050d0402", 
1422 => x"f0050d75", 
1423 => x"5372802e", 
1424 => x"a13872bd", 
1425 => x"980c80c1", 
1426 => x"bc08fe14", 
1427 => x"712980c1", 
1428 => x"c0080580", 
1429 => x"c1b40c70", 
1430 => x"842b80c1", 
1431 => x"a00c54ad", 
1432 => x"8e04bd9c", 
1433 => x"08bd980c", 
1434 => x"80c1a808", 
1435 => x"80c1b40c", 
1436 => x"80c1b008", 
1437 => x"802e8b38", 
1438 => x"80c1bc08", 
1439 => x"842b53ad", 
1440 => x"890480c1", 
1441 => x"b808842b", 
1442 => x"537280c1", 
1443 => x"a00c0290", 
1444 => x"050d0402", 
1445 => x"ec050d76", 
1446 => x"5574802e", 
1447 => x"80e93874", 
1448 => x"84e02d54", 
1449 => x"73802e80", 
1450 => x"de389ce0", 
1451 => x"528151a3", 
1452 => x"8f2d8808", 
1453 => x"54880880", 
1454 => x"2e80cc38", 
1455 => x"8b537452", 
1456 => x"8808519c", 
1457 => x"a32d8808", 
1458 => x"802e8938", 
1459 => x"9ce05280", 
1460 => x"51adaf04", 
1461 => x"73802eaf", 
1462 => x"389a1480", 
1463 => x"c02d5194", 
1464 => x"c42d8808", 
1465 => x"5580c1b0", 
1466 => x"08802e96", 
1467 => x"38941480", 
1468 => x"c02d5194", 
1469 => x"c42d8808", 
1470 => x"902b83ff", 
1471 => x"f00a0675", 
1472 => x"05557451", 
1473 => x"acb72d02", 
1474 => x"94050d04", 
1475 => x"02f8050d", 
1476 => x"bd980870", 
1477 => x"535170bd", 
1478 => x"9c082e09", 
1479 => x"81068338", 
1480 => x"80527188", 
1481 => x"0c028805", 
1482 => x"0d0402f4", 
1483 => x"050d7452", 
1484 => x"80537173", 
1485 => x"2eaa389a", 
1486 => x"1280c02d", 
1487 => x"5194c42d", 
1488 => x"88085380", 
1489 => x"c1b00880", 
1490 => x"2e963894", 
1491 => x"1280c02d", 
1492 => x"5194c42d", 
1493 => x"8808902b", 
1494 => x"83fff00a", 
1495 => x"06730753", 
1496 => x"7251acb7", 
1497 => x"2d028c05", 
1498 => x"0d0402e8", 
1499 => x"050d7856", 
1500 => x"80785255", 
1501 => x"acb72daf", 
1502 => x"b2048808", 
1503 => x"9a0580c0", 
1504 => x"2d5194c4", 
1505 => x"2d880854", 
1506 => x"80c1b008", 
1507 => x"802e9638", 
1508 => x"941580c0", 
1509 => x"2d5194c4", 
1510 => x"2d880890", 
1511 => x"2b83fff0", 
1512 => x"0a067405", 
1513 => x"5473762e", 
1514 => x"09810686", 
1515 => x"388153af", 
1516 => x"cd048052", 
1517 => x"74810509", 
1518 => x"70760780", 
1519 => x"255253a3", 
1520 => x"8f2d8808", 
1521 => x"558808ff", 
1522 => x"b1388808", 
1523 => x"5372880c", 
1524 => x"0298050d", 
1525 => x"0402d805", 
1526 => x"0d7b5978", 
1527 => x"802e8b38", 
1528 => x"78bd9c08", 
1529 => x"2e098106", 
1530 => x"86388154", 
1531 => x"b1b504fe", 
1532 => x"1980c1bc", 
1533 => x"082980c1", 
1534 => x"c00811bd", 
1535 => x"a0545254", 
1536 => x"93c62d88", 
1537 => x"08548808", 
1538 => x"802e81a9", 
1539 => x"38bda056", 
1540 => x"80588076", 
1541 => x"84e02d55", 
1542 => x"5573752e", 
1543 => x"83388155", 
1544 => x"7381e52e", 
1545 => x"81813881", 
1546 => x"70760655", 
1547 => x"5a73802e", 
1548 => x"80f5388b", 
1549 => x"1684e02d", 
1550 => x"70842a70", 
1551 => x"7c065155", 
1552 => x"5573802e", 
1553 => x"80e13888", 
1554 => x"53b8a852", 
1555 => x"7551b3a5", 
1556 => x"2d880857", 
1557 => x"880880cf", 
1558 => x"389a1680", 
1559 => x"c02d5194", 
1560 => x"c42d8808", 
1561 => x"88085555", 
1562 => x"80c1b008", 
1563 => x"802e9738", 
1564 => x"941680c0", 
1565 => x"2d5194c4", 
1566 => x"2d880890", 
1567 => x"2b83fff0", 
1568 => x"0a067016", 
1569 => x"51547674", 
1570 => x"5255afd5", 
1571 => x"2d880880", 
1572 => x"2e903878", 
1573 => x"527351ae", 
1574 => x"ea2d8808", 
1575 => x"802e8338", 
1576 => x"79557454", 
1577 => x"b1b504a0", 
1578 => x"16811959", 
1579 => x"568f7827", 
1580 => x"fee03880", 
1581 => x"5473880c", 
1582 => x"02a8050d", 
1583 => x"04fb3d0d", 
1584 => x"77795555", 
1585 => x"80567476", 
1586 => x"25863874", 
1587 => x"30558156", 
1588 => x"73802588", 
1589 => x"38733076", 
1590 => x"81325754", 
1591 => x"80537352", 
1592 => x"745180ca", 
1593 => x"3f880854", 
1594 => x"75802e85", 
1595 => x"38880830", 
1596 => x"5473880c", 
1597 => x"873d0d04", 
1598 => x"fa3d0d78", 
1599 => x"7a575580", 
1600 => x"57747725", 
1601 => x"86387430", 
1602 => x"55815775", 
1603 => x"9f2c5481", 
1604 => x"53757432", 
1605 => x"74315274", 
1606 => x"51943f88", 
1607 => x"08547680", 
1608 => x"2e853888", 
1609 => x"08305473", 
1610 => x"880c883d", 
1611 => x"0d04fc3d", 
1612 => x"0d767853", 
1613 => x"54815380", 
1614 => x"55873971", 
1615 => x"10731054", 
1616 => x"52737226", 
1617 => x"5172802e", 
1618 => x"a7387080", 
1619 => x"2e863871", 
1620 => x"8025e838", 
1621 => x"72802e98", 
1622 => x"38717426", 
1623 => x"89387372", 
1624 => x"31757407", 
1625 => x"56547281", 
1626 => x"2a72812a", 
1627 => x"5353e539", 
1628 => x"73517883", 
1629 => x"38745170", 
1630 => x"880c863d", 
1631 => x"0d04fd3d", 
1632 => x"0d757754", 
1633 => x"52805471", 
1634 => x"8106ff11", 
1635 => x"70097506", 
1636 => x"1674812a", 
1637 => x"76105755", 
1638 => x"56515171", 
1639 => x"ea387388", 
1640 => x"0c853d0d", 
1641 => x"04fc3d0d", 
1642 => x"76787a70", 
1643 => x"55535454", 
1644 => x"70802eb6", 
1645 => x"389f3973", 
1646 => x"33733356", 
1647 => x"5271752e", 
1648 => x"0981069c", 
1649 => x"3870802e", 
1650 => x"97387180", 
1651 => x"2e923881", 
1652 => x"14811454", 
1653 => x"54ff1151", 
1654 => x"70ff2e09", 
1655 => x"8106d838", 
1656 => x"73337333", 
1657 => x"71713154", 
1658 => x"54547188", 
1659 => x"0c863d0d", 
1660 => x"04fe3d0d", 
1661 => x"74b58511", 
1662 => x"3370812a", 
1663 => x"70810651", 
1664 => x"53545270", 
1665 => x"802e8438", 
1666 => x"e0125271", 
1667 => x"880c843d", 
1668 => x"0d040000", 
1669 => x"00ffffff", 
1670 => x"ff00ffff", 
1671 => x"ffff00ff", 
1672 => x"ffffff00", 
1673 => x"4f4e4452", 
1674 => x"41202020", 
1675 => x"20202000", 
1676 => x"00000000", 
1677 => x"00000bbd", 
1678 => x"00000b73", 
1679 => x"00000be2", 
1680 => x"00000c56", 
1681 => x"00000d47", 
1682 => x"00000d5e", 
1683 => x"00000b73", 
1684 => x"00000b73", 
1685 => x"00000db2", 
1686 => x"00000b73", 
1687 => x"00000dd7", 
1688 => x"00000ddc", 
1689 => x"00000de1", 
1690 => x"00000dec", 
1691 => x"00000b73", 
1692 => x"00000df1", 
1693 => x"00000b73", 
1694 => x"00000b73", 
1695 => x"00000b73", 
1696 => x"00000df6", 
1697 => x"00202020", 
1698 => x"20202020", 
1699 => x"20202828", 
1700 => x"28282820", 
1701 => x"20202020", 
1702 => x"20202020", 
1703 => x"20202020", 
1704 => x"20202020", 
1705 => x"20881010", 
1706 => x"10101010", 
1707 => x"10101010", 
1708 => x"10101010", 
1709 => x"10040404", 
1710 => x"04040404", 
1711 => x"04040410", 
1712 => x"10101010", 
1713 => x"10104141", 
1714 => x"41414141", 
1715 => x"01010101", 
1716 => x"01010101", 
1717 => x"01010101", 
1718 => x"01010101", 
1719 => x"01010101", 
1720 => x"10101010", 
1721 => x"10104242", 
1722 => x"42424242", 
1723 => x"02020202", 
1724 => x"02020202", 
1725 => x"02020202", 
1726 => x"02020202", 
1727 => x"02020202", 
1728 => x"10101010", 
1729 => x"20000000", 
1730 => x"00000000", 
1731 => x"00000000", 
1732 => x"00000000", 
1733 => x"00000000", 
1734 => x"00000000", 
1735 => x"00000000", 
1736 => x"00000000", 
1737 => x"00000000", 
1738 => x"00000000", 
1739 => x"00000000", 
1740 => x"00000000", 
1741 => x"00000000", 
1742 => x"00000000", 
1743 => x"00000000", 
1744 => x"00000000", 
1745 => x"00000000", 
1746 => x"00000000", 
1747 => x"00000000", 
1748 => x"00000000", 
1749 => x"00000000", 
1750 => x"00000000", 
1751 => x"00000000", 
1752 => x"00000000", 
1753 => x"00000000", 
1754 => x"00000000", 
1755 => x"00000000", 
1756 => x"00000000", 
1757 => x"00000000", 
1758 => x"00000000", 
1759 => x"00000000", 
1760 => x"00000000", 
1761 => x"00000000", 
1762 => x"5f5f4c4f", 
1763 => x"41444552", 
1764 => x"42494e00", 
1765 => x"2f202020", 
1766 => x"20202020", 
1767 => x"20202000", 
1768 => x"2e202020", 
1769 => x"20202020", 
1770 => x"20202000", 
1771 => x"54415000", 
1772 => x"0a0d4f6e", 
1773 => x"64726153", 
1774 => x"4420696e", 
1775 => x"74657266", 
1776 => x"61636520", 
1777 => x"28322e32", 
1778 => x"29202b20", 
1779 => x"5254430a", 
1780 => x"0d4d3120", 
1781 => x"28632920", 
1782 => x"32303135", 
1783 => x"2c203230", 
1784 => x"31360a0d", 
1785 => x"68747470", 
1786 => x"733a2f2f", 
1787 => x"73697465", 
1788 => x"732e676f", 
1789 => x"6f676c65", 
1790 => x"2e636f6d", 
1791 => x"2f736974", 
1792 => x"652f6f6e", 
1793 => x"64726173", 
1794 => x"706f3138", 
1795 => x"360a0d00", 
1796 => x"46415431", 
1797 => x"36202020", 
1798 => x"00000000", 
1799 => x"46415433", 
1800 => x"32202020", 
1801 => x"00000000", 
1802 => x"2e2e2020", 
1803 => x"20202020", 
1804 => x"20202000", 
1805 => x"000000fa", 
1806 => x"00001c10", 
1807 => x"00001c1c", 
1808 => x"ffffffff", 
1809 => x"00001a85", 


	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

