-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity Ondra_TESLA_V5 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(11 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of Ondra_TESLA_V5 is


  type ROM_ARRAY is array(0 to 4095) of std_logic_vector(7 downto 0);
  constant ROM : ROM_ARRAY := (
    x"F3",x"AF",x"D3",x"03",x"C3",x"CB",x"24",x"00", -- 0x0000
    x"C3",x"AE",x"00",x"32",x"4D",x"03",x"C9",x"00", -- 0x0008
    x"E3",x"7E",x"E6",x"7F",x"CD",x"B3",x"05",x"7E", -- 0x0010
    x"07",x"23",x"30",x"F5",x"E3",x"C9",x"3E",x"01", -- 0x0018
    x"FB",x"E5",x"21",x"B8",x"CE",x"86",x"BE",x"20", -- 0x0020
    x"FD",x"E1",x"C9",x"AF",x"B9",x"3E",x"02",x"28", -- 0x0028
    x"03",x"3E",x"03",x"FB",x"D3",x"03",x"C9",x"00", -- 0x0030
    x"08",x"D9",x"3E",x"07",x"D3",x"03",x"01",x"0A", -- 0x0038
    x"00",x"11",x"A9",x"CE",x"21",x"00",x"E0",x"ED", -- 0x0040
    x"B0",x"3E",x"03",x"D3",x"03",x"D9",x"3A",x"B8", -- 0x0048
    x"CE",x"3C",x"32",x"B8",x"CE",x"08",x"FB",x"C9", -- 0x0050
    x"21",x"7F",x"CE",x"AF",x"77",x"23",x"BD",x"20", -- 0x0058
    x"FB",x"21",x"7F",x"CE",x"18",x"02",x"18",x"07", -- 0x0060
    x"22",x"D9",x"CE",x"F9",x"CD",x"93",x"01",x"21", -- 0x0068
    x"80",x"CE",x"22",x"A0",x"CE",x"D7",x"0D",x"0A", -- 0x0070
    x"4F",x"6E",x"64",x"72",x"61",x"20",x"56",x"2E", -- 0x0078
    x"35",x"87",x"AF",x"32",x"CC",x"CE",x"31",x"94", -- 0x0080
    x"CE",x"AF",x"32",x"A2",x"CE",x"3D",x"32",x"A7", -- 0x0088
    x"CE",x"CD",x"C3",x"06",x"21",x"AE",x"00",x"22", -- 0x0090
    x"09",x"00",x"21",x"86",x"00",x"E5",x"CD",x"C8", -- 0x0098
    x"03",x"D7",x"0D",x"0A",x"AE",x"CD",x"3A",x"06", -- 0x00A0
    x"FE",x"43",x"C2",x"16",x"05",x"C7",x"F3",x"22", -- 0x00A8
    x"9C",x"CE",x"EB",x"22",x"9A",x"CE",x"F5",x"21", -- 0x00B0
    x"02",x"00",x"39",x"22",x"A0",x"CE",x"F1",x"E1", -- 0x00B8
    x"22",x"9E",x"CE",x"31",x"9A",x"CE",x"C5",x"F5", -- 0x00C0
    x"CD",x"77",x"05",x"18",x"B9",x"21",x"DB",x"CE", -- 0x00C8
    x"11",x"D1",x"CE",x"06",x"06",x"1A",x"4E",x"77", -- 0x00D0
    x"79",x"12",x"23",x"13",x"10",x"F7",x"C9",x"CD", -- 0x00D8
    x"F0",x"05",x"CD",x"14",x"06",x"D7",x"A0",x"C9", -- 0x00E0
    x"CD",x"E6",x"08",x"CD",x"1E",x"00",x"3A",x"AC", -- 0x00E8
    x"CE",x"E6",x"40",x"20",x"F3",x"79",x"D3",x"09", -- 0x00F0
    x"AF",x"D3",x"0A",x"C3",x"ED",x"01",x"00",x"00", -- 0x00F8
    x"C7",x"64",x"04",x"C3",x"16",x"03",x"C3",x"20", -- 0x0100
    x"0A",x"C3",x"9B",x"01",x"C3",x"6B",x"0A",x"C3", -- 0x0108
    x"EB",x"00",x"C3",x"46",x"03",x"C3",x"6A",x"06", -- 0x0110
    x"C3",x"31",x"00",x"C3",x"52",x"06",x"C3",x"5A", -- 0x0118
    x"06",x"C3",x"63",x"06",x"C3",x"F0",x"05",x"C3", -- 0x0120
    x"CB",x"05",x"C3",x"AA",x"05",x"C3",x"27",x"06", -- 0x0128
    x"C3",x"E2",x"00",x"C3",x"19",x"06",x"C3",x"FB", -- 0x0130
    x"05",x"C3",x"86",x"00",x"C3",x"E5",x"00",x"C3", -- 0x0138
    x"3A",x"06",x"C3",x"49",x"06",x"C3",x"19",x"05", -- 0x0140
    x"C3",x"0C",x"06",x"C3",x"6E",x"06",x"C3",x"E2", -- 0x0148
    x"01",x"C3",x"2B",x"00",x"C3",x"77",x"09",x"C3", -- 0x0150
    x"69",x"07",x"C3",x"9D",x"0C",x"C3",x"06",x"0C", -- 0x0158
    x"C3",x"5F",x"0C",x"C3",x"D0",x"00",x"3E",x"42", -- 0x0160
    x"32",x"E4",x"CE",x"C9",x"7C",x"BA",x"CC",x"79", -- 0x0168
    x"01",x"C8",x"3D",x"16",x"7A",x"32",x"D2",x"CE", -- 0x0170
    x"C9",x"7D",x"BB",x"C8",x"B7",x"C8",x"3D",x"32", -- 0x0178
    x"D1",x"CE",x"3A",x"D6",x"CE",x"B7",x"C0",x"3E", -- 0x0180
    x"28",x"B7",x"C9",x"CD",x"74",x"01",x"7B",x"32", -- 0x0188
    x"D1",x"CE",x"C9",x"21",x"E7",x"FF",x"22",x"A3", -- 0x0190
    x"CE",x"0E",x"1F",x"E5",x"D5",x"C5",x"21",x"AD", -- 0x0198
    x"02",x"E5",x"2A",x"A3",x"CE",x"3A",x"A5",x"CE", -- 0x01A0
    x"77",x"79",x"FE",x"20",x"30",x"49",x"2A",x"D3", -- 0x01A8
    x"CE",x"EB",x"2A",x"D1",x"CE",x"FE",x"0D",x"28", -- 0x01B0
    x"BB",x"FE",x"0A",x"28",x"53",x"FE",x"1E",x"CA", -- 0x01B8
    x"55",x"02",x"FE",x"08",x"28",x"A6",x"FE",x"1D", -- 0x01C0
    x"28",x"C1",x"FE",x"1F",x"CA",x"6A",x"02",x"FE", -- 0x01C8
    x"18",x"28",x"2A",x"FE",x"1A",x"28",x"A2",x"FE", -- 0x01D0
    x"1C",x"CA",x"CD",x"00",x"FE",x"07",x"C0",x"01", -- 0x01D8
    x"05",x"05",x"78",x"0F",x"0F",x"0F",x"E6",x"E0", -- 0x01E0
    x"CD",x"F2",x"01",x"79",x"E7",x"3A",x"A2",x"CE", -- 0x01E8
    x"E6",x"03",x"F6",x"08",x"D3",x"0A",x"C9",x"CD", -- 0x01F0
    x"CF",x"02",x"CD",x"FB",x"02",x"2A",x"D1",x"CE", -- 0x01F8
    x"24",x"22",x"D1",x"CE",x"CD",x"82",x"01",x"3D", -- 0x0200
    x"BC",x"D0",x"3A",x"D4",x"CE",x"32",x"D2",x"CE", -- 0x0208
    x"CD",x"96",x"02",x"47",x"7D",x"3C",x"B8",x"DA", -- 0x0210
    x"8F",x"01",x"2A",x"D3",x"CE",x"E5",x"CD",x"96", -- 0x0218
    x"02",x"47",x"3E",x"18",x"90",x"85",x"6F",x"CD", -- 0x0220
    x"ED",x"02",x"0F",x"D6",x"80",x"4F",x"E1",x"CD", -- 0x0228
    x"ED",x"02",x"0F",x"D6",x"80",x"6F",x"CD",x"9E", -- 0x0230
    x"02",x"06",x"00",x"C5",x"F5",x"E5",x"C5",x"CD", -- 0x0238
    x"7B",x"02",x"C1",x"E1",x"E5",x"3E",x"80",x"85", -- 0x0240
    x"6F",x"03",x"CD",x"7B",x"02",x"E1",x"F1",x"C1", -- 0x0248
    x"25",x"BC",x"20",x"E7",x"C9",x"CD",x"ED",x"02", -- 0x0250
    x"CD",x"9E",x"02",x"BC",x"C8",x"F5",x"E5",x"11", -- 0x0258
    x"00",x"D0",x"CD",x"FB",x"02",x"E1",x"F1",x"25", -- 0x0260
    x"18",x"F1",x"E5",x"CD",x"55",x"02",x"E1",x"3A", -- 0x0268
    x"D4",x"CE",x"67",x"CD",x"96",x"02",x"2C",x"BD", -- 0x0270
    x"20",x"F0",x"C9",x"54",x"3E",x"05",x"85",x"5F", -- 0x0278
    x"ED",x"B8",x"CD",x"8C",x"02",x"06",x"06",x"71", -- 0x0280
    x"23",x"10",x"FC",x"C9",x"01",x"00",x"0A",x"3A", -- 0x0288
    x"CC",x"CE",x"07",x"D0",x"0D",x"C9",x"3A",x"D5", -- 0x0290
    x"CE",x"B7",x"C0",x"3E",x"18",x"C9",x"E5",x"CD", -- 0x0298
    x"82",x"01",x"67",x"CD",x"ED",x"02",x"7C",x"E1", -- 0x02A0
    x"FE",x"D7",x"C0",x"3D",x"C9",x"3A",x"CC",x"CE", -- 0x02A8
    x"0F",x"C1",x"C5",x"F5",x"DC",x"0F",x"01",x"CD", -- 0x02B0
    x"EA",x"02",x"CB",x"0D",x"22",x"A3",x"CE",x"7E", -- 0x02B8
    x"32",x"A5",x"CE",x"F1",x"0F",x"38",x"03",x"7E", -- 0x02C0
    x"2F",x"77",x"C1",x"D1",x"E1",x"79",x"C9",x"79", -- 0x02C8
    x"11",x"00",x"D0",x"D6",x"21",x"38",x"13",x"3C", -- 0x02D0
    x"26",x"00",x"F2",x"DF",x"02",x"D6",x"40",x"D5", -- 0x02D8
    x"6F",x"29",x"54",x"5D",x"29",x"29",x"19",x"D1", -- 0x02E0
    x"19",x"EB",x"2A",x"D1",x"CE",x"7C",x"2F",x"67", -- 0x02E8
    x"7D",x"07",x"47",x"07",x"07",x"80",x"2F",x"C6", -- 0x02F0
    x"E8",x"6F",x"C9",x"CD",x"8C",x"02",x"CB",x"0D", -- 0x02F8
    x"1A",x"A9",x"77",x"13",x"CB",x"05",x"2C",x"10", -- 0x0300
    x"F5",x"C9",x"3A",x"CC",x"CE",x"A8",x"32",x"CC", -- 0x0308
    x"CE",x"C1",x"3C",x"CC",x"AE",x"00",x"FB",x"C5", -- 0x0310
    x"D5",x"E5",x"CD",x"4C",x"03",x"E1",x"D1",x"78", -- 0x0318
    x"06",x"01",x"FE",x"10",x"28",x"E4",x"06",x"80", -- 0x0320
    x"FE",x"12",x"28",x"DE",x"C1",x"FE",x"17",x"28", -- 0x0328
    x"E2",x"FE",x"11",x"C0",x"CD",x"16",x"03",x"FE", -- 0x0330
    x"47",x"20",x"04",x"3E",x"16",x"18",x"02",x"E6", -- 0x0338
    x"0F",x"32",x"D3",x"CE",x"18",x"D0",x"E5",x"CD", -- 0x0340
    x"CB",x"03",x"E1",x"C9",x"0E",x"01",x"CD",x"CB", -- 0x0348
    x"03",x"20",x"02",x"0E",x"08",x"CD",x"C8",x"03", -- 0x0350
    x"EB",x"C4",x"C8",x"03",x"28",x"F5",x"CD",x"00", -- 0x0358
    x"06",x"20",x"F0",x"44",x"7D",x"D6",x"A9",x"6F", -- 0x0360
    x"87",x"87",x"85",x"5F",x"16",x"00",x"D5",x"21", -- 0x0368
    x"34",x"04",x"3A",x"A2",x"CE",x"E6",x"03",x"87", -- 0x0370
    x"5F",x"19",x"5E",x"23",x"56",x"EB",x"D1",x"19", -- 0x0378
    x"78",x"06",x"05",x"0F",x"30",x"05",x"2B",x"10", -- 0x0380
    x"FA",x"18",x"C8",x"79",x"3D",x"C4",x"20",x"00", -- 0x0388
    x"3A",x"A2",x"CE",x"F5",x"01",x"01",x"01",x"CD", -- 0x0390
    x"E2",x"01",x"32",x"A2",x"CE",x"F1",x"FE",x"04", -- 0x0398
    x"20",x"10",x"7E",x"E6",x"3F",x"47",x"FE",x"0D", -- 0x03A0
    x"20",x"02",x"06",x"1D",x"FE",x"0A",x"C0",x"06", -- 0x03A8
    x"1F",x"C9",x"46",x"0F",x"30",x"0A",x"F5",x"3E", -- 0x03B0
    x"40",x"B8",x"30",x"03",x"0F",x"80",x"47",x"F1", -- 0x03B8
    x"E6",x"40",x"C8",x"78",x"EE",x"A0",x"47",x"C9", -- 0x03C0
    x"CD",x"1E",x"00",x"D5",x"C5",x"21",x"AD",x"CE", -- 0x03C8
    x"7E",x"F6",x"E9",x"2E",x"AB",x"CB",x"66",x"20", -- 0x03D0
    x"02",x"E6",x"F7",x"2E",x"B0",x"CB",x"66",x"20", -- 0x03D8
    x"01",x"3D",x"21",x"A7",x"CE",x"46",x"77",x"B8", -- 0x03E0
    x"30",x"08",x"A8",x"CD",x"0D",x"04",x"77",x"CD", -- 0x03E8
    x"ED",x"01",x"11",x"A9",x"CE",x"21",x"D2",x"04", -- 0x03F0
    x"1A",x"A6",x"BE",x"20",x"06",x"23",x"13",x"7E", -- 0x03F8
    x"3C",x"20",x"F5",x"67",x"6B",x"C4",x"ED",x"01", -- 0x0400
    x"C1",x"D1",x"7C",x"B7",x"C9",x"21",x"A2",x"CE", -- 0x0408
    x"0F",x"30",x"03",x"3E",x"04",x"C9",x"0F",x"30", -- 0x0410
    x"09",x"7E",x"E6",x"03",x"D6",x"03",x"C8",x"3E", -- 0x0418
    x"03",x"C9",x"0F",x"30",x"06",x"7E",x"E6",x"FD", -- 0x0420
    x"F6",x"80",x"C9",x"0F",x"06",x"02",x"38",x"01", -- 0x0428
    x"05",x"7E",x"A8",x"C9",x"40",x"04",x"40",x"04", -- 0x0430
    x"72",x"04",x"A4",x"04",x"51",x"54",x"57",x"45", -- 0x0438
    x"52",x"41",x"47",x"53",x"44",x"46",x"00",x"56", -- 0x0440
    x"5A",x"58",x"43",x"00",x"00",x"00",x"00",x"20", -- 0x0448
    x"00",x"00",x"00",x"00",x"00",x"0D",x"48",x"4C", -- 0x0450
    x"4B",x"4A",x"50",x"59",x"4F",x"49",x"55",x"00", -- 0x0458
    x"42",x"1A",x"4D",x"4E",x"18",x"00",x"0A",x"08", -- 0x0460
    x"00",x"0D",x"0A",x"1A",x"08",x"18",x"21",x"25", -- 0x0468
    x"22",x"23",x"24",x"2D",x"5F",x"2B",x"3D",x"5E", -- 0x0470
    x"00",x"3B",x"2A",x"2F",x"3A",x"00",x"00",x"00", -- 0x0478
    x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"0D", -- 0x0480
    x"3C",x"5D",x"5B",x"3E",x"40",x"26",x"29",x"28", -- 0x0488
    x"27",x"00",x"3F",x"1A",x"2E",x"2C",x"18",x"00", -- 0x0490
    x"0A",x"08",x"00",x"0D",x"0A",x"1A",x"08",x"18", -- 0x0498
    x"31",x"35",x"32",x"33",x"34",x"2D",x"5F",x"2B", -- 0x04A0
    x"3D",x"5E",x"00",x"3B",x"2A",x"2F",x"3A",x"00", -- 0x04A8
    x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00", -- 0x04B0
    x"00",x"0D",x"3C",x"5D",x"5B",x"3E",x"30",x"36", -- 0x04B8
    x"39",x"38",x"37",x"00",x"3F",x"1A",x"2E",x"2C", -- 0x04C0
    x"18",x"00",x"0A",x"08",x"00",x"0D",x"0A",x"1A", -- 0x04C8
    x"08",x"18",x"1F",x"1F",x"0F",x"03",x"00",x"1F", -- 0x04D0
    x"1F",x"0F",x"1F",x"1F",x"FF",x"0E",x"03",x"CD", -- 0x04D8
    x"CB",x"05",x"C1",x"D1",x"E1",x"7E",x"02",x"03", -- 0x04E0
    x"CD",x"FB",x"05",x"30",x"F8",x"C9",x"CD",x"BA", -- 0x04E8
    x"05",x"7D",x"E6",x"07",x"CC",x"DF",x"00",x"7E", -- 0x04F0
    x"CD",x"19",x"06",x"CD",x"38",x"06",x"D8",x"28", -- 0x04F8
    x"0D",x"FE",x"08",x"2B",x"28",x"EE",x"23",x"EB", -- 0x0500
    x"CD",x"C1",x"05",x"EB",x"73",x"C8",x"23",x"FE", -- 0x0508
    x"2C",x"CC",x"DF",x"00",x"18",x"DB",x"2A",x"9E", -- 0x0510
    x"CE",x"FE",x"4D",x"28",x"C0",x"FE",x"47",x"28", -- 0x0518
    x"2F",x"FE",x"53",x"28",x"C9",x"FE",x"58",x"28", -- 0x0520
    x"49",x"FE",x"4B",x"CA",x"7F",x"06",x"FE",x"4C", -- 0x0528
    x"CA",x"F7",x"0B",x"FE",x"42",x"C2",x"84",x"06", -- 0x0530
    x"2A",x"B3",x"CE",x"7E",x"FE",x"C3",x"C2",x"6F", -- 0x0538
    x"00",x"3A",x"A8",x"CE",x"B7",x"20",x"05",x"3D", -- 0x0540
    x"32",x"A8",x"CE",x"E9",x"23",x"23",x"23",x"E9", -- 0x0548
    x"CD",x"BA",x"05",x"22",x"9E",x"CE",x"CD",x"F0", -- 0x0550
    x"05",x"31",x"96",x"CE",x"F1",x"C1",x"D1",x"2A", -- 0x0558
    x"A0",x"CE",x"F9",x"2A",x"9E",x"CE",x"E3",x"2A", -- 0x0560
    x"9C",x"CE",x"C9",x"41",x"42",x"44",x"48",x"50", -- 0x0568
    x"53",x"00",x"CD",x"3A",x"06",x"30",x"04",x"CD", -- 0x0570
    x"F0",x"05",x"3E",x"AF",x"32",x"A6",x"CE",x"11", -- 0x0578
    x"96",x"CE",x"01",x"6B",x"05",x"0A",x"B7",x"C8", -- 0x0580
    x"CD",x"B3",x"05",x"D7",x"AD",x"03",x"1A",x"6F", -- 0x0588
    x"13",x"1A",x"67",x"C5",x"D7",x"A0",x"CD",x"E2", -- 0x0590
    x"00",x"3A",x"A6",x"CE",x"B7",x"CC",x"BD",x"05", -- 0x0598
    x"C1",x"1B",x"7D",x"12",x"13",x"7C",x"12",x"13", -- 0x05A0
    x"18",x"DB",x"D7",x"07",x"BF",x"C3",x"6F",x"00", -- 0x05A8
    x"CD",x"16",x"03",x"C5",x"4F",x"CD",x"9B",x"01", -- 0x05B0
    x"C1",x"C9",x"CD",x"E2",x"00",x"CD",x"38",x"06", -- 0x05B8
    x"C8",x"CD",x"F4",x"05",x"E1",x"78",x"FE",x"0D", -- 0x05C0
    x"C9",x"38",x"DF",x"D7",x"BD",x"21",x"00",x"00", -- 0x05C8
    x"CD",x"B0",x"05",x"47",x"CD",x"27",x"06",x"38", -- 0x05D0
    x"0B",x"29",x"29",x"29",x"29",x"B5",x"6F",x"3E", -- 0x05D8
    x"02",x"E7",x"18",x"EC",x"78",x"CD",x"3D",x"06", -- 0x05E0
    x"20",x"C0",x"E3",x"E5",x"0D",x"20",x"DA",x"D0", -- 0x05E8
    x"D7",x"0D",x"8A",x"C9",x"0E",x"01",x"21",x"00", -- 0x05F0
    x"00",x"18",x"D8",x"23",x"7C",x"B5",x"37",x"C8", -- 0x05F8
    x"7A",x"BC",x"C0",x"7B",x"BD",x"C9",x"0F",x"0F", -- 0x0600
    x"0F",x"0F",x"E6",x"0F",x"C6",x"90",x"27",x"CE", -- 0x0608
    x"40",x"27",x"4F",x"C9",x"7C",x"CD",x"19",x"06", -- 0x0610
    x"7D",x"F5",x"CD",x"06",x"06",x"CD",x"9B",x"01", -- 0x0618
    x"F1",x"CD",x"0A",x"06",x"C3",x"9B",x"01",x"D6", -- 0x0620
    x"30",x"D8",x"FE",x"17",x"3F",x"D8",x"FE",x"0A", -- 0x0628
    x"3F",x"D0",x"FE",x"11",x"D8",x"D6",x"07",x"C9", -- 0x0630
    x"D7",x"AD",x"CD",x"B0",x"05",x"FE",x"2C",x"C8", -- 0x0638
    x"FE",x"20",x"C8",x"FE",x"0D",x"37",x"C8",x"B7", -- 0x0640
    x"C9",x"4E",x"23",x"CD",x"9B",x"01",x"15",x"20", -- 0x0648
    x"F8",x"C9",x"E5",x"2A",x"D9",x"CE",x"7D",x"44", -- 0x0650
    x"E1",x"C9",x"3E",x"08",x"B9",x"C0",x"EB",x"22", -- 0x0658
    x"D9",x"CE",x"C9",x"2A",x"D1",x"CE",x"EB",x"2A", -- 0x0660
    x"A3",x"CE",x"3A",x"D3",x"CE",x"C9",x"47",x"79", -- 0x0668
    x"FE",x"0C",x"78",x"D0",x"E5",x"06",x"00",x"21", -- 0x0670
    x"CC",x"CE",x"09",x"77",x"EB",x"E1",x"C9",x"D7", -- 0x0678
    x"DF",x"CD",x"30",x"09",x"F5",x"3E",x"14",x"E7", -- 0x0680
    x"F1",x"32",x"D7",x"CE",x"FE",x"41",x"CA",x"79", -- 0x0688
    x"07",x"FE",x"44",x"28",x"49",x"FE",x"49",x"CA", -- 0x0690
    x"4B",x"08",x"FE",x"4F",x"28",x"64",x"FE",x"43", -- 0x0698
    x"CA",x"9D",x"0C",x"FE",x"46",x"CA",x"7C",x"09", -- 0x06A0
    x"FE",x"53",x"CA",x"5F",x"0C",x"FE",x"4C",x"CA", -- 0x06A8
    x"06",x"0C",x"FE",x"4A",x"28",x"23",x"FE",x"54", -- 0x06B0
    x"28",x"12",x"FE",x"4D",x"C0",x"CD",x"0D",x"09", -- 0x06B8
    x"CD",x"22",x"09",x"C5",x"CD",x"31",x"00",x"CD", -- 0x06C0
    x"ED",x"01",x"C1",x"C9",x"2A",x"B3",x"CE",x"CD", -- 0x06C8
    x"DF",x"00",x"EB",x"2A",x"B5",x"CE",x"C3",x"E2", -- 0x06D0
    x"00",x"CD",x"CC",x"06",x"EB",x"E9",x"CD",x"01", -- 0x06D8
    x"09",x"3C",x"CC",x"CF",x"08",x"AF",x"2A",x"EF", -- 0x06E0
    x"CF",x"22",x"C5",x"CE",x"0E",x"24",x"C4",x"09", -- 0x06E8
    x"01",x"CD",x"39",x"09",x"28",x"EC",x"FE",x"04", -- 0x06F0
    x"D5",x"CC",x"2A",x"08",x"D1",x"CD",x"17",x"0A", -- 0x06F8
    x"18",x"E4",x"AF",x"32",x"D7",x"CE",x"3A",x"CF", -- 0x0700
    x"CE",x"B7",x"20",x"76",x"CD",x"8F",x"07",x"28", -- 0x0708
    x"0C",x"D7",x"0D",x"0A",x"70",x"6F",x"73",x"6C", -- 0x0710
    x"65",x"64",x"6E",x"69",x"A0",x"CD",x"95",x"07", -- 0x0718
    x"20",x"14",x"CD",x"39",x"09",x"28",x"0C",x"FE", -- 0x0720
    x"04",x"20",x"F7",x"CD",x"1E",x"08",x"CD",x"39", -- 0x0728
    x"08",x"28",x"14",x"CD",x"E3",x"07",x"C4",x"E0", -- 0x0730
    x"07",x"3A",x"E4",x"CE",x"FE",x"3A",x"28",x"07", -- 0x0738
    x"CD",x"39",x"09",x"FE",x"04",x"20",x"F9",x"7A", -- 0x0740
    x"3C",x"67",x"2E",x"00",x"22",x"C5",x"CE",x"CD", -- 0x0748
    x"1A",x"09",x"CD",x"8F",x"07",x"28",x"07",x"D7", -- 0x0750
    x"0D",x"0A",x"6E",x"6F",x"76",x"F9",x"3E",x"01", -- 0x0758
    x"32",x"CF",x"CE",x"32",x"E4",x"CE",x"C3",x"7A", -- 0x0760
    x"08",x"CD",x"87",x"07",x"FE",x"22",x"20",x"96", -- 0x0768
    x"23",x"7E",x"FE",x"40",x"20",x"90",x"22",x"C9", -- 0x0770
    x"CE",x"32",x"B9",x"CE",x"2A",x"C5",x"CE",x"EB", -- 0x0778
    x"18",x"C5",x"CD",x"9D",x"0C",x"18",x"F2",x"7E", -- 0x0780
    x"32",x"D7",x"CE",x"22",x"C9",x"CE",x"C9",x"3A", -- 0x0788
    x"D7",x"CE",x"FE",x"22",x"C9",x"3E",x"AF",x"32", -- 0x0790
    x"B9",x"CE",x"B7",x"F5",x"CD",x"8F",x"07",x"F5", -- 0x0798
    x"C4",x"DC",x"08",x"21",x"BA",x"CE",x"06",x"0B", -- 0x07A0
    x"F1",x"20",x"08",x"F1",x"36",x"2A",x"CC",x"C4", -- 0x07A8
    x"07",x"18",x"04",x"CD",x"AD",x"08",x"F1",x"CD", -- 0x07B0
    x"01",x"09",x"21",x"BA",x"CE",x"7E",x"FE",x"2A", -- 0x07B8
    x"C8",x"FE",x"0D",x"C9",x"D5",x"EB",x"2A",x"C9", -- 0x07C0
    x"CE",x"EB",x"13",x"1A",x"77",x"B7",x"28",x"09", -- 0x07C8
    x"FE",x"22",x"28",x"05",x"23",x"10",x"F3",x"D1", -- 0x07D0
    x"C9",x"36",x"20",x"D1",x"C9",x"CD",x"CF",x"08", -- 0x07D8
    x"CD",x"39",x"09",x"20",x"FB",x"FE",x"3A",x"20", -- 0x07E0
    x"06",x"3A",x"B9",x"CE",x"B7",x"28",x"EE",x"01", -- 0x07E8
    x"BA",x"CE",x"1E",x"0B",x"23",x"0A",x"FE",x"2A", -- 0x07F0
    x"28",x"19",x"CD",x"40",x"06",x"28",x"07",x"BE", -- 0x07F8
    x"20",x"DE",x"03",x"1D",x"20",x"EE",x"D5",x"D7", -- 0x0800
    x"87",x"21",x"E4",x"CE",x"E5",x"CD",x"CF",x"08", -- 0x0808
    x"E1",x"D1",x"C9",x"CD",x"06",x"08",x"CD",x"39", -- 0x0810
    x"08",x"20",x"C5",x"C9",x"D7",x"9D",x"21",x"E4", -- 0x0818
    x"CF",x"16",x"0B",x"CD",x"49",x"06",x"2A",x"EF", -- 0x0820
    x"CF",x"EB",x"D7",x"A0",x"7A",x"CD",x"19",x"06", -- 0x0828
    x"D7",x"AD",x"7B",x"CD",x"19",x"06",x"D7",x"9E", -- 0x0830
    x"C9",x"D7",x"07",x"2D",x"2D",x"28",x"59",x"2F", -- 0x0838
    x"4E",x"29",x"BF",x"CD",x"30",x"09",x"E6",x"DF", -- 0x0840
    x"FE",x"59",x"C9",x"CD",x"0D",x"09",x"D7",x"70", -- 0x0848
    x"72",x"65",x"76",x"69",x"6E",x"20",x"2D",x"20", -- 0x0850
    x"7A",x"61",x"70",x"6E",x"69",x"A0",x"CD",x"1A", -- 0x0858
    x"09",x"CD",x"C3",x"06",x"D7",x"20",x"7A",x"61", -- 0x0860
    x"64",x"65",x"6A",x"A0",x"21",x"00",x"00",x"22", -- 0x0868
    x"C5",x"CE",x"3E",x"3A",x"32",x"E4",x"CE",x"32", -- 0x0870
    x"D7",x"CE",x"CD",x"8F",x"07",x"F5",x"C4",x"DC", -- 0x0878
    x"08",x"CD",x"0A",x"0A",x"CD",x"C3",x"06",x"23", -- 0x0880
    x"06",x"40",x"F1",x"E5",x"F5",x"C4",x"AD",x"08", -- 0x0888
    x"F1",x"CC",x"C4",x"07",x"E1",x"06",x"0B",x"11", -- 0x0890
    x"F4",x"CF",x"7E",x"E6",x"7F",x"20",x"02",x"3E", -- 0x0898
    x"20",x"12",x"23",x"13",x"10",x"F4",x"CD",x"FF", -- 0x08A0
    x"09",x"36",x"41",x"18",x"1F",x"5D",x"D7",x"BA", -- 0x08A8
    x"36",x"20",x"CD",x"EF",x"08",x"FE",x"0D",x"28", -- 0x08B0
    x"13",x"FE",x"08",x"20",x"0B",x"7B",x"BD",x"28", -- 0x08B8
    x"ED",x"2B",x"04",x"D7",x"20",x"88",x"18",x"E8", -- 0x08C0
    x"77",x"23",x"10",x"E4",x"C3",x"F0",x"05",x"CD", -- 0x08C8
    x"F0",x"05",x"23",x"16",x"40",x"CD",x"49",x"06", -- 0x08D0
    x"3E",x"64",x"E7",x"C9",x"D7",x"20",x"6E",x"61", -- 0x08D8
    x"7A",x"65",x"76",x"0D",x"8A",x"C9",x"CD",x"46", -- 0x08E0
    x"03",x"C8",x"CD",x"03",x"01",x"18",x"04",x"CD", -- 0x08E8
    x"3A",x"06",x"C8",x"F5",x"3E",x"02",x"E7",x"F1", -- 0x08F0
    x"FE",x"03",x"C0",x"CD",x"4F",x"0C",x"C3",x"86", -- 0x08F8
    x"00",x"D7",x"20",x"63",x"74",x"65",x"6E",x"69", -- 0x0900
    x"20",x"AD",x"CD",x"22",x"09",x"3A",x"CB",x"CE", -- 0x0908
    x"B7",x"3E",x"19",x"28",x"02",x"3E",x"1B",x"D3", -- 0x0910
    x"0A",x"C9",x"D7",x"20",x"7A",x"61",x"70",x"69", -- 0x0918
    x"73",x"A1",x"D7",x"20",x"68",x"6F",x"74",x"6F", -- 0x0920
    x"76",x"6F",x"BF",x"CD",x"46",x"03",x"28",x"FB", -- 0x0928
    x"CD",x"EF",x"08",x"F5",x"CD",x"F0",x"05",x"F1", -- 0x0930
    x"C9",x"AF",x"0E",x"23",x"DC",x"09",x"01",x"CD", -- 0x0938
    x"6F",x"09",x"CD",x"62",x"0B",x"F5",x"E5",x"21", -- 0x0940
    x"CC",x"CE",x"7E",x"F5",x"36",x"80",x"2A",x"D1", -- 0x0948
    x"CE",x"E5",x"CD",x"31",x"00",x"CD",x"1C",x"08", -- 0x0950
    x"E1",x"22",x"D1",x"CE",x"F1",x"32",x"CC",x"CE", -- 0x0958
    x"3A",x"B7",x"CE",x"B7",x"C4",x"EF",x"08",x"20", -- 0x0960
    x"FB",x"E1",x"F1",x"38",x"CD",x"18",x"37",x"2A", -- 0x0968
    x"C5",x"CE",x"23",x"22",x"C5",x"CE",x"C9",x"CD", -- 0x0970
    x"87",x"07",x"18",x"04",x"AF",x"32",x"D7",x"CE", -- 0x0978
    x"CD",x"96",x"07",x"CD",x"E0",x"07",x"1E",x"01", -- 0x0980
    x"EB",x"22",x"C5",x"CE",x"EB",x"3E",x"01",x"32", -- 0x0988
    x"B9",x"CE",x"32",x"CD",x"CE",x"D5",x"C5",x"CD", -- 0x0990
    x"6F",x"09",x"CD",x"66",x"0B",x"38",x"0F",x"CD", -- 0x0998
    x"17",x"0A",x"20",x"0A",x"C1",x"D1",x"7E",x"FE", -- 0x09A0
    x"3A",x"C8",x"FE",x"01",x"C9",x"F1",x"CD",x"C3", -- 0x09A8
    x"06",x"2A",x"C5",x"CE",x"CD",x"DF",x"00",x"D7", -- 0x09B0
    x"0D",x"0A",x"07",x"43",x"68",x"79",x"62",x"61", -- 0x09B8
    x"20",x"63",x"74",x"65",x"6E",x"69",x"20",x"2D", -- 0x09C0
    x"20",x"5A",x"6E",x"6F",x"76",x"61",x"2F",x"4E", -- 0x09C8
    x"BF",x"CD",x"EF",x"08",x"E6",x"DF",x"FE",x"4E", -- 0x09D0
    x"28",x"20",x"D7",x"20",x"76",x"72",x"61",x"74", -- 0x09D8
    x"20",x"7A",x"70",x"65",x"74",x"A0",x"CD",x"01", -- 0x09E0
    x"09",x"CD",x"62",x"0B",x"F5",x"CD",x"17",x"0A", -- 0x09E8
    x"28",x"05",x"30",x"B9",x"F1",x"18",x"F2",x"F1", -- 0x09F0
    x"38",x"B4",x"CD",x"F0",x"05",x"18",x"A5",x"D5", -- 0x09F8
    x"C5",x"CD",x"6F",x"09",x"EB",x"CD",x"8B",x"0A", -- 0x0A00
    x"C1",x"D1",x"21",x"E4",x"CE",x"E5",x"06",x"FF", -- 0x0A08
    x"23",x"36",x"00",x"10",x"FB",x"E1",x"C9",x"E5", -- 0x0A10
    x"2A",x"C5",x"CE",x"CD",x"00",x"06",x"E1",x"C9", -- 0x0A18
    x"C5",x"D5",x"E5",x"3A",x"CD",x"CE",x"B7",x"CC", -- 0x0A20
    x"7C",x"09",x"2A",x"C7",x"CE",x"23",x"7D",x"FE", -- 0x0A28
    x"E4",x"7E",x"22",x"C7",x"CE",x"28",x"1F",x"FE", -- 0x0A30
    x"1A",x"20",x"2B",x"4F",x"CD",x"50",x"0A",x"79", -- 0x0A38
    x"20",x"24",x"5D",x"21",x"E4",x"CF",x"2B",x"BE", -- 0x0A40
    x"20",x"FC",x"7D",x"93",x"20",x"F1",x"18",x"0F", -- 0x0A48
    x"3A",x"E4",x"CE",x"FE",x"04",x"C9",x"CD",x"50", -- 0x0A50
    x"0A",x"C4",x"95",x"09",x"20",x"CF",x"AF",x"32", -- 0x0A58
    x"CD",x"CE",x"3E",x"1A",x"37",x"06",x"B7",x"E1", -- 0x0A60
    x"D1",x"C1",x"C9",x"C5",x"D5",x"E5",x"3A",x"CF", -- 0x0A68
    x"CE",x"B7",x"C5",x"CC",x"02",x"07",x"C1",x"2A", -- 0x0A70
    x"C7",x"CE",x"23",x"71",x"22",x"C7",x"CE",x"7D", -- 0x0A78
    x"FE",x"E3",x"CC",x"FF",x"09",x"E1",x"D1",x"C1", -- 0x0A80
    x"79",x"B7",x"C9",x"EB",x"22",x"EF",x"CF",x"21", -- 0x0A88
    x"F4",x"CF",x"11",x"E4",x"CF",x"01",x"0B",x"00", -- 0x0A90
    x"ED",x"B0",x"CD",x"E6",x"08",x"21",x"10",x"10", -- 0x0A98
    x"22",x"E1",x"CE",x"22",x"E2",x"CE",x"22",x"F2", -- 0x0AA0
    x"CF",x"CD",x"4D",x"0B",x"78",x"32",x"F1",x"CF", -- 0x0AA8
    x"21",x"E1",x"CE",x"CD",x"15",x"09",x"3A",x"E4", -- 0x0AB0
    x"CE",x"FE",x"3A",x"20",x"08",x"F5",x"3E",x"FF", -- 0x0AB8
    x"E7",x"3E",x"FF",x"E7",x"F1",x"FE",x"42",x"28", -- 0x0AC0
    x"03",x"3E",x"28",x"E7",x"F3",x"11",x"C2",x"03", -- 0x0AC8
    x"01",x"13",x"01",x"3E",x"06",x"D3",x"03",x"3E", -- 0x0AD0
    x"01",x"CD",x"31",x"0B",x"1B",x"7B",x"B2",x"20", -- 0x0AD8
    x"F6",x"7E",x"23",x"CD",x"16",x"0B",x"0B",x"79", -- 0x0AE0
    x"B0",x"20",x"F6",x"01",x"0A",x"00",x"11",x"A9", -- 0x0AE8
    x"CE",x"21",x"00",x"E0",x"ED",x"B0",x"2A",x"EF", -- 0x0AF0
    x"CF",x"EB",x"21",x"E4",x"CE",x"22",x"C7",x"CE", -- 0x0AF8
    x"7E",x"FE",x"42",x"F5",x"3E",x"0B",x"20",x"02", -- 0x0B00
    x"3E",x"18",x"D3",x"0A",x"7E",x"FE",x"04",x"CC", -- 0x0B08
    x"ED",x"01",x"F1",x"C3",x"2D",x"00",x"C5",x"F5", -- 0x0B10
    x"4F",x"AF",x"CD",x"31",x"0B",x"06",x"08",x"79", -- 0x0B18
    x"CD",x"31",x"0B",x"0F",x"10",x"FA",x"3E",x"01", -- 0x0B20
    x"CD",x"31",x"0B",x"CD",x"31",x"0B",x"F1",x"C1", -- 0x0B28
    x"C9",x"C5",x"F5",x"07",x"07",x"07",x"E6",x"08", -- 0x0B30
    x"F6",x"02",x"D3",x"03",x"EE",x"08",x"0E",x"19", -- 0x0B38
    x"0D",x"20",x"FD",x"D3",x"03",x"0E",x"11",x"0D", -- 0x0B40
    x"20",x"FD",x"F1",x"C1",x"C9",x"D5",x"21",x"E4", -- 0x0B48
    x"CE",x"01",x"0D",x"01",x"16",x"00",x"7A",x"86", -- 0x0B50
    x"57",x"23",x"0B",x"78",x"B1",x"20",x"F7",x"42", -- 0x0B58
    x"D1",x"C9",x"AF",x"32",x"CB",x"CE",x"C5",x"21", -- 0x0B60
    x"E4",x"CE",x"CD",x"0D",x"09",x"3E",x"06",x"D3", -- 0x0B68
    x"03",x"F3",x"06",x"1E",x"CD",x"D8",x"0B",x"38", -- 0x0B70
    x"F9",x"10",x"F9",x"06",x"03",x"CD",x"BD",x"0B", -- 0x0B78
    x"FE",x"10",x"20",x"EE",x"10",x"F7",x"01",x"0F", -- 0x0B80
    x"01",x"CD",x"BD",x"0B",x"77",x"23",x"0B",x"79", -- 0x0B88
    x"B0",x"20",x"F6",x"CD",x"EB",x"0A",x"E5",x"3A", -- 0x0B90
    x"F2",x"CF",x"FE",x"10",x"20",x"17",x"CD",x"E6", -- 0x0B98
    x"08",x"28",x"01",x"3E",x"AF",x"32",x"B7",x"CE", -- 0x0BA0
    x"3D",x"32",x"CB",x"CE",x"CD",x"4D",x"0B",x"3A", -- 0x0BA8
    x"F1",x"CF",x"90",x"28",x"01",x"37",x"2A",x"EF", -- 0x0BB0
    x"CF",x"EB",x"E1",x"C1",x"C9",x"C5",x"06",x"80", -- 0x0BB8
    x"CD",x"D8",x"0B",x"30",x"FB",x"4F",x"CD",x"D8", -- 0x0BC0
    x"0B",x"D4",x"D8",x"0B",x"A9",x"07",x"CB",x"18", -- 0x0BC8
    x"30",x"F4",x"CD",x"D8",x"0B",x"78",x"C1",x"C9", -- 0x0BD0
    x"E5",x"C5",x"06",x"0E",x"21",x"03",x"E0",x"4E", -- 0x0BD8
    x"7E",x"A9",x"F2",x"E8",x"0B",x"A9",x"18",x"0A", -- 0x0BE0
    x"05",x"20",x"F5",x"7E",x"A9",x"F2",x"EB",x"0B", -- 0x0BE8
    x"A9",x"37",x"C1",x"E1",x"C9",x"22",x"0D",x"21", -- 0x0BF0
    x"F5",x"0B",x"AF",x"32",x"A8",x"CE",x"CD",x"06", -- 0x0BF8
    x"0C",x"3E",x"42",x"C3",x"38",x"05",x"CD",x"77", -- 0x0C00
    x"09",x"CD",x"0D",x"09",x"23",x"7E",x"D6",x"3C", -- 0x0C08
    x"20",x"47",x"2A",x"E6",x"CE",x"22",x"B5",x"CE", -- 0x0C10
    x"E5",x"2A",x"E8",x"CE",x"22",x"B3",x"CE",x"3E", -- 0x0C18
    x"0D",x"94",x"30",x"35",x"EB",x"3A",x"EA",x"CE", -- 0x0C20
    x"FE",x"3E",x"20",x"2D",x"01",x"F8",x"00",x"21", -- 0x0C28
    x"EC",x"CE",x"CD",x"50",x"0A",x"28",x"0C",x"ED", -- 0x0C30
    x"B0",x"CD",x"95",x"09",x"21",x"E5",x"CE",x"0E", -- 0x0C38
    x"FF",x"18",x"EF",x"44",x"4D",x"EB",x"D1",x"0A", -- 0x0C40
    x"77",x"03",x"CD",x"FB",x"05",x"30",x"F8",x"AF", -- 0x0C48
    x"32",x"CD",x"CE",x"CD",x"C3",x"06",x"C3",x"F0", -- 0x0C50
    x"05",x"CD",x"4F",x"0C",x"C3",x"AA",x"05",x"0E", -- 0x0C58
    x"02",x"CD",x"CB",x"05",x"3A",x"CF",x"CE",x"B7", -- 0x0C60
    x"CC",x"02",x"07",x"CD",x"66",x"01",x"CD",x"0D", -- 0x0C68
    x"09",x"3E",x"28",x"E7",x"0E",x"3C",x"CD",x"C5", -- 0x0C70
    x"0C",x"06",x"00",x"E1",x"D1",x"CD",x"C0",x"0C", -- 0x0C78
    x"EB",x"CD",x"C0",x"0C",x"0E",x"3E",x"CD",x"C5", -- 0x0C80
    x"0C",x"48",x"CD",x"C5",x"0C",x"06",x"00",x"4E", -- 0x0C88
    x"CD",x"C5",x"0C",x"CD",x"FB",x"05",x"D2",x"8F", -- 0x0C90
    x"0C",x"48",x"CD",x"C5",x"0C",x"3A",x"CF",x"CE", -- 0x0C98
    x"B7",x"CA",x"AA",x"05",x"E5",x"0E",x"1A",x"CD", -- 0x0CA0
    x"6B",x"0A",x"3E",x"04",x"32",x"E4",x"CE",x"CD", -- 0x0CA8
    x"FF",x"09",x"AF",x"32",x"CF",x"CE",x"CD",x"0D", -- 0x0CB0
    x"09",x"3E",x"28",x"E7",x"E1",x"C3",x"C3",x"06", -- 0x0CB8
    x"4D",x"CD",x"C5",x"0C",x"4C",x"79",x"80",x"47", -- 0x0CC0
    x"C3",x"6B",x"0A",x"3C",x"D3",x"0A",x"3E",x"30", -- 0x0CC8
    x"D3",x"03",x"3E",x"14",x"DB",x"09",x"3E",x"7A", -- 0x0CD0
    x"DB",x"3D",x"3E",x"B2",x"DB",x"5A",x"AF",x"D3", -- 0x0CD8
    x"03",x"3E",x"40",x"DB",x"78",x"3E",x"10",x"D3", -- 0x0CE0
    x"03",x"3E",x"2F",x"DB",x"06",x"AF",x"DB",x"80", -- 0x0CE8
    x"3E",x"20",x"D3",x"03",x"3E",x"29",x"DB",x"1C", -- 0x0CF0
    x"AF",x"DB",x"80",x"21",x"00",x"D0",x"AF",x"77", -- 0x0CF8
    x"23",x"BC",x"20",x"FB",x"3E",x"3E",x"21",x"4E", -- 0x0D00
    x"25",x"11",x"0B",x"D0",x"01",x"07",x"00",x"ED", -- 0x0D08
    x"B0",x"13",x"13",x"13",x"3D",x"20",x"F5",x"3D", -- 0x0D10
    x"12",x"11",x"80",x"D2",x"21",x"00",x"27",x"3E", -- 0x0D18
    x"20",x"01",x"08",x"00",x"ED",x"B0",x"13",x"13", -- 0x0D20
    x"3D",x"20",x"F6",x"11",x"00",x"80",x"63",x"6B", -- 0x0D28
    x"01",x"00",x"08",x"ED",x"B0",x"44",x"26",x"20", -- 0x0D30
    x"ED",x"B0",x"C3",x"3D",x"8D",x"3E",x"02",x"D3", -- 0x0D38
    x"03",x"53",x"26",x"80",x"01",x"CB",x"0C",x"ED", -- 0x0D40
    x"B0",x"ED",x"56",x"C3",x"58",x"00",x"30",x"00", -- 0x0D48
    x"30",x"30",x"78",x"78",x"30",x"00",x"00",x"00", -- 0x0D50
    x"00",x"6C",x"6C",x"6C",x"6C",x"6C",x"FE",x"6C", -- 0x0D58
    x"FE",x"6C",x"6C",x"30",x"F8",x"0C",x"78",x"C0", -- 0x0D60
    x"7C",x"30",x"C6",x"66",x"30",x"18",x"CC",x"C6", -- 0x0D68
    x"00",x"76",x"CC",x"DC",x"76",x"38",x"6C",x"38", -- 0x0D70
    x"00",x"00",x"00",x"00",x"C0",x"60",x"60",x"18", -- 0x0D78
    x"30",x"60",x"60",x"60",x"30",x"18",x"60",x"30", -- 0x0D80
    x"18",x"18",x"18",x"30",x"60",x"00",x"66",x"3C", -- 0x0D88
    x"FF",x"3C",x"66",x"00",x"00",x"30",x"30",x"FC", -- 0x0D90
    x"30",x"30",x"00",x"60",x"30",x"30",x"00",x"00", -- 0x0D98
    x"00",x"00",x"00",x"00",x"00",x"FC",x"00",x"00", -- 0x0DA0
    x"00",x"30",x"30",x"00",x"00",x"00",x"00",x"00", -- 0x0DA8
    x"80",x"C0",x"60",x"30",x"18",x"0C",x"06",x"7C", -- 0x0DB0
    x"E6",x"F6",x"DE",x"CE",x"C6",x"7C",x"FC",x"30", -- 0x0DB8
    x"30",x"30",x"30",x"70",x"30",x"FC",x"CC",x"60", -- 0x0DC0
    x"38",x"0C",x"CC",x"78",x"78",x"CC",x"0C",x"38", -- 0x0DC8
    x"0C",x"CC",x"78",x"1E",x"0C",x"FE",x"CC",x"6C", -- 0x0DD0
    x"3C",x"1C",x"78",x"CC",x"0C",x"0C",x"F8",x"C0", -- 0x0DD8
    x"FC",x"78",x"CC",x"CC",x"F8",x"C0",x"60",x"38", -- 0x0DE0
    x"30",x"30",x"30",x"18",x"0C",x"CC",x"FC",x"78", -- 0x0DE8
    x"CC",x"CC",x"78",x"CC",x"CC",x"78",x"70",x"18", -- 0x0DF0
    x"0C",x"7C",x"CC",x"CC",x"78",x"30",x"30",x"00", -- 0x0DF8
    x"00",x"30",x"30",x"00",x"60",x"30",x"30",x"00", -- 0x0E00
    x"30",x"30",x"00",x"18",x"30",x"60",x"C0",x"60", -- 0x0E08
    x"30",x"18",x"00",x"FC",x"00",x"00",x"FC",x"00", -- 0x0E10
    x"00",x"60",x"30",x"18",x"0C",x"18",x"30",x"60", -- 0x0E18
    x"30",x"00",x"30",x"18",x"0C",x"CC",x"78",x"78", -- 0x0E20
    x"C0",x"DE",x"DE",x"DE",x"C6",x"7C",x"CC",x"CC", -- 0x0E28
    x"FC",x"CC",x"CC",x"78",x"30",x"FC",x"66",x"66", -- 0x0E30
    x"7C",x"66",x"66",x"FC",x"3C",x"66",x"C0",x"C0", -- 0x0E38
    x"C0",x"66",x"3C",x"F8",x"6C",x"66",x"66",x"66", -- 0x0E40
    x"6C",x"F8",x"FE",x"62",x"68",x"78",x"68",x"62", -- 0x0E48
    x"FE",x"F0",x"60",x"68",x"78",x"68",x"62",x"FE", -- 0x0E50
    x"3E",x"66",x"CE",x"C0",x"C0",x"66",x"3C",x"CC", -- 0x0E58
    x"CC",x"CC",x"FC",x"CC",x"CC",x"CC",x"78",x"30", -- 0x0E60
    x"30",x"30",x"30",x"30",x"78",x"78",x"CC",x"CC", -- 0x0E68
    x"0C",x"0C",x"0C",x"1E",x"E6",x"66",x"6C",x"78", -- 0x0E70
    x"6C",x"66",x"E6",x"FE",x"66",x"62",x"60",x"60", -- 0x0E78
    x"60",x"F0",x"C6",x"C6",x"D6",x"FE",x"FE",x"EE", -- 0x0E80
    x"C6",x"C6",x"C6",x"CE",x"DE",x"F6",x"E6",x"C6", -- 0x0E88
    x"38",x"6C",x"C6",x"C6",x"C6",x"6C",x"38",x"F0", -- 0x0E90
    x"60",x"60",x"7C",x"66",x"66",x"FC",x"1C",x"78", -- 0x0E98
    x"DC",x"CC",x"CC",x"CC",x"78",x"E6",x"66",x"6C", -- 0x0EA0
    x"7C",x"66",x"66",x"FC",x"78",x"CC",x"1C",x"70", -- 0x0EA8
    x"E0",x"CC",x"78",x"78",x"30",x"30",x"30",x"30", -- 0x0EB0
    x"B4",x"FC",x"FC",x"CC",x"CC",x"CC",x"CC",x"CC", -- 0x0EB8
    x"CC",x"30",x"78",x"CC",x"CC",x"CC",x"CC",x"CC", -- 0x0EC0
    x"C6",x"EE",x"FE",x"D6",x"C6",x"C6",x"C6",x"C6", -- 0x0EC8
    x"6C",x"38",x"38",x"6C",x"C6",x"C6",x"78",x"30", -- 0x0ED0
    x"30",x"78",x"CC",x"CC",x"CC",x"FE",x"66",x"32", -- 0x0ED8
    x"18",x"8C",x"C6",x"FE",x"78",x"60",x"60",x"60", -- 0x0EE0
    x"60",x"60",x"78",x"02",x"06",x"0C",x"18",x"30", -- 0x0EE8
    x"60",x"C0",x"78",x"18",x"18",x"18",x"18",x"18", -- 0x0EF0
    x"78",x"00",x"00",x"00",x"C6",x"6C",x"38",x"10", -- 0x0EF8
    x"00",x"00",x"00",x"00",x"00",x"18",x"30",x"30", -- 0x0F00
    x"00",x"76",x"CC",x"7C",x"0C",x"78",x"00",x"00", -- 0x0F08
    x"00",x"DC",x"66",x"66",x"7C",x"60",x"60",x"E0", -- 0x0F10
    x"00",x"78",x"CC",x"C0",x"CC",x"78",x"00",x"00", -- 0x0F18
    x"00",x"76",x"CC",x"CC",x"7C",x"0C",x"0C",x"1C", -- 0x0F20
    x"00",x"78",x"C0",x"FC",x"CC",x"78",x"00",x"00", -- 0x0F28
    x"00",x"F0",x"60",x"60",x"F0",x"60",x"6C",x"38", -- 0x0F30
    x"F8",x"0C",x"7C",x"CC",x"CC",x"76",x"00",x"00", -- 0x0F38
    x"00",x"E6",x"66",x"66",x"76",x"6C",x"60",x"E0", -- 0x0F40
    x"00",x"78",x"30",x"30",x"30",x"70",x"00",x"30", -- 0x0F48
    x"78",x"CC",x"CC",x"0C",x"0C",x"0C",x"00",x"0C", -- 0x0F50
    x"00",x"E6",x"6C",x"78",x"6C",x"66",x"60",x"E0", -- 0x0F58
    x"00",x"78",x"30",x"30",x"30",x"30",x"30",x"70", -- 0x0F60
    x"00",x"C6",x"D6",x"FE",x"FE",x"CC",x"00",x"00", -- 0x0F68
    x"00",x"CC",x"CC",x"CC",x"CC",x"F8",x"00",x"00", -- 0x0F70
    x"00",x"78",x"CC",x"CC",x"CC",x"78",x"00",x"00", -- 0x0F78
    x"F0",x"60",x"7C",x"66",x"66",x"DC",x"00",x"00", -- 0x0F80
    x"1E",x"0C",x"7C",x"CC",x"CC",x"76",x"00",x"00", -- 0x0F88
    x"00",x"F0",x"60",x"66",x"76",x"DC",x"00",x"00", -- 0x0F90
    x"00",x"F8",x"0C",x"78",x"C0",x"7C",x"00",x"00", -- 0x0F98
    x"00",x"18",x"34",x"30",x"30",x"7C",x"30",x"10", -- 0x0FA0
    x"00",x"76",x"CC",x"CC",x"CC",x"CC",x"00",x"00", -- 0x0FA8
    x"00",x"30",x"78",x"CC",x"CC",x"CC",x"00",x"00", -- 0x0FB0
    x"00",x"6C",x"FE",x"FE",x"D6",x"C6",x"00",x"00", -- 0x0FB8
    x"00",x"C6",x"6C",x"38",x"6C",x"C6",x"00",x"00", -- 0x0FC0
    x"F8",x"0C",x"7C",x"CC",x"CC",x"CC",x"00",x"00", -- 0x0FC8
    x"00",x"FC",x"64",x"30",x"98",x"FC",x"00",x"00", -- 0x0FD0
    x"00",x"1C",x"30",x"30",x"E0",x"30",x"30",x"1C", -- 0x0FD8
    x"00",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0FE0
    x"00",x"E0",x"30",x"30",x"1C",x"30",x"30",x"E0", -- 0x0FE8
    x"00",x"00",x"00",x"00",x"00",x"00",x"DC",x"76", -- 0x0FF0
    x"00",x"FE",x"C6",x"C6",x"6C",x"38",x"10",x"00"  -- 0x0FF8
  );

begin

  p_rom : process
  begin
    wait until rising_edge(CLK);
    if (ENA = '1') then
       DATA <= ROM(to_integer(unsigned(ADDR)));
    end if;
  end process;
end RTL;
